/* ============================================================================
 *  Title       : Prime number ROM
 *
 *  File Name	: PRIME_ROM.v
 *  Project     :
 *  Block       :
 *  Tree        :
 *  Designer    : toms74209200 <https://github.com/toms74209200>
 *  Created     : 2019/09/22
 *  Copyright   : 2019 toms74209200
 *  License     : MIT License.
 *                http://opensource.org/licenses/mit-license.php
 * ============================================================================*/
module PRIME_ROM
    (
    // System
    CLK,        //(p) Clock

    // ROM interface
    ADDRESS,    //(p) Address
    DATA        //(p) Data
    );

// Port
// System
input           CLK;        //(p) Clock

// ROM interface
input  [10:0]   ADDRESS;    //(p) Address
output [15:0]   DATA;       //(p) Data

// Internal signals
reg [15:0]      data_i;     // Data

/* ============================================================================
 * ROM output
 * ============================================================================*/
always@(posedge CLK) begin
    case (ADDRESS)
        0   : data_i <= 16'h0003;
        1   : data_i <= 16'h0005;
        2   : data_i <= 16'h0007;
        3   : data_i <= 16'h000B;
        4   : data_i <= 16'h000D;
        5   : data_i <= 16'h0011;
        6   : data_i <= 16'h0013;
        7   : data_i <= 16'h0017;
        8   : data_i <= 16'h001D;
        9   : data_i <= 16'h001F;
        10  : data_i <= 16'h0025;
        11  : data_i <= 16'h0029;
        12  : data_i <= 16'h002B;
        13  : data_i <= 16'h002F;
        14  : data_i <= 16'h0035;
        15  : data_i <= 16'h003B;
        16  : data_i <= 16'h003D;
        17  : data_i <= 16'h0043;
        18  : data_i <= 16'h0047;
        19  : data_i <= 16'h0049;
        20  : data_i <= 16'h004F;
        21  : data_i <= 16'h0053;
        22  : data_i <= 16'h0059;
        23  : data_i <= 16'h0061;
        24  : data_i <= 16'h0065;
        25  : data_i <= 16'h0067;
        26  : data_i <= 16'h006B;
        27  : data_i <= 16'h006D;
        28  : data_i <= 16'h0071;
        29  : data_i <= 16'h007F;
        30  : data_i <= 16'h0083;
        31  : data_i <= 16'h0089;
        32  : data_i <= 16'h008B;
        33  : data_i <= 16'h0095;
        34  : data_i <= 16'h0097;
        35  : data_i <= 16'h009D;
        36  : data_i <= 16'h00A3;
        37  : data_i <= 16'h00A7;
        38  : data_i <= 16'h00AD;
        39  : data_i <= 16'h00B3;
        40  : data_i <= 16'h00B5;
        41  : data_i <= 16'h00BF;
        42  : data_i <= 16'h00C1;
        43  : data_i <= 16'h00C5;
        44  : data_i <= 16'h00C7;
        45  : data_i <= 16'h00D3;
        46  : data_i <= 16'h00DF;
        47  : data_i <= 16'h00E3;
        48  : data_i <= 16'h00E5;
        49  : data_i <= 16'h00E9;
        50  : data_i <= 16'h00EF;
        51  : data_i <= 16'h00F1;
        52  : data_i <= 16'h00FB;
        53  : data_i <= 16'h0101;
        54  : data_i <= 16'h0107;
        55  : data_i <= 16'h010D;
        56  : data_i <= 16'h010F;
        57  : data_i <= 16'h0115;
        58  : data_i <= 16'h0119;
        59  : data_i <= 16'h011B;
        60  : data_i <= 16'h0125;
        61  : data_i <= 16'h0133;
        62  : data_i <= 16'h0137;
        63  : data_i <= 16'h0139;
        64  : data_i <= 16'h013D;
        65  : data_i <= 16'h014B;
        66  : data_i <= 16'h0151;
        67  : data_i <= 16'h015B;
        68  : data_i <= 16'h015D;
        69  : data_i <= 16'h0161;
        70  : data_i <= 16'h0167;
        71  : data_i <= 16'h016F;
        72  : data_i <= 16'h0175;
        73  : data_i <= 16'h017B;
        74  : data_i <= 16'h017F;
        75  : data_i <= 16'h0185;
        76  : data_i <= 16'h018D;
        77  : data_i <= 16'h0191;
        78  : data_i <= 16'h0199;
        79  : data_i <= 16'h01A3;
        80  : data_i <= 16'h01A5;
        81  : data_i <= 16'h01AF;
        82  : data_i <= 16'h01B1;
        83  : data_i <= 16'h01B7;
        84  : data_i <= 16'h01BB;
        85  : data_i <= 16'h01C1;
        86  : data_i <= 16'h01C9;
        87  : data_i <= 16'h01CD;
        88  : data_i <= 16'h01CF;
        89  : data_i <= 16'h01D3;
        90  : data_i <= 16'h01DF;
        91  : data_i <= 16'h01E7;
        92  : data_i <= 16'h01EB;
        93  : data_i <= 16'h01F3;
        94  : data_i <= 16'h01F7;
        95  : data_i <= 16'h01FD;
        96  : data_i <= 16'h0209;
        97  : data_i <= 16'h020B;
        98  : data_i <= 16'h021D;
        99  : data_i <= 16'h0223;
        100 : data_i <= 16'h022D;
        101 : data_i <= 16'h0233;
        102 : data_i <= 16'h0239;
        103 : data_i <= 16'h023B;
        104 : data_i <= 16'h0241;
        105 : data_i <= 16'h024B;
        106 : data_i <= 16'h0251;
        107 : data_i <= 16'h0257;
        108 : data_i <= 16'h0259;
        109 : data_i <= 16'h025F;
        110 : data_i <= 16'h0265;
        111 : data_i <= 16'h0269;
        112 : data_i <= 16'h026B;
        113 : data_i <= 16'h0277;
        114 : data_i <= 16'h0281;
        115 : data_i <= 16'h0283;
        116 : data_i <= 16'h0287;
        117 : data_i <= 16'h028D;
        118 : data_i <= 16'h0293;
        119 : data_i <= 16'h0295;
        120 : data_i <= 16'h02A1;
        121 : data_i <= 16'h02A5;
        122 : data_i <= 16'h02AB;
        123 : data_i <= 16'h02B3;
        124 : data_i <= 16'h02BD;
        125 : data_i <= 16'h02C5;
        126 : data_i <= 16'h02CF;
        127 : data_i <= 16'h02D7;
        128 : data_i <= 16'h02DD;
        129 : data_i <= 16'h02E3;
        130 : data_i <= 16'h02E7;
        131 : data_i <= 16'h02EF;
        132 : data_i <= 16'h02F5;
        133 : data_i <= 16'h02F9;
        134 : data_i <= 16'h0301;
        135 : data_i <= 16'h0305;
        136 : data_i <= 16'h0313;
        137 : data_i <= 16'h031D;
        138 : data_i <= 16'h0329;
        139 : data_i <= 16'h032B;
        140 : data_i <= 16'h0335;
        141 : data_i <= 16'h0337;
        142 : data_i <= 16'h033B;
        143 : data_i <= 16'h033D;
        144 : data_i <= 16'h0347;
        145 : data_i <= 16'h0355;
        146 : data_i <= 16'h0359;
        147 : data_i <= 16'h035B;
        148 : data_i <= 16'h035F;
        149 : data_i <= 16'h036D;
        150 : data_i <= 16'h0371;
        151 : data_i <= 16'h0373;
        152 : data_i <= 16'h0377;
        153 : data_i <= 16'h038B;
        154 : data_i <= 16'h038F;
        155 : data_i <= 16'h0397;
        156 : data_i <= 16'h03A1;
        157 : data_i <= 16'h03A9;
        158 : data_i <= 16'h03AD;
        159 : data_i <= 16'h03B3;
        160 : data_i <= 16'h03B9;
        161 : data_i <= 16'h03C7;
        162 : data_i <= 16'h03CB;
        163 : data_i <= 16'h03D1;
        164 : data_i <= 16'h03D7;
        165 : data_i <= 16'h03DF;
        166 : data_i <= 16'h03E5;
        167 : data_i <= 16'h03F1;
        168 : data_i <= 16'h03F5;
        169 : data_i <= 16'h03FB;
        170 : data_i <= 16'h03FD;
        171 : data_i <= 16'h0407;
        172 : data_i <= 16'h0409;
        173 : data_i <= 16'h040F;
        174 : data_i <= 16'h0419;
        175 : data_i <= 16'h041B;
        176 : data_i <= 16'h0425;
        177 : data_i <= 16'h0427;
        178 : data_i <= 16'h042D;
        179 : data_i <= 16'h043F;
        180 : data_i <= 16'h0443;
        181 : data_i <= 16'h0445;
        182 : data_i <= 16'h0449;
        183 : data_i <= 16'h044F;
        184 : data_i <= 16'h0455;
        185 : data_i <= 16'h045D;
        186 : data_i <= 16'h0463;
        187 : data_i <= 16'h0469;
        188 : data_i <= 16'h047F;
        189 : data_i <= 16'h0481;
        190 : data_i <= 16'h048B;
        191 : data_i <= 16'h0493;
        192 : data_i <= 16'h049D;
        193 : data_i <= 16'h04A3;
        194 : data_i <= 16'h04A9;
        195 : data_i <= 16'h04B1;
        196 : data_i <= 16'h04BD;
        197 : data_i <= 16'h04C1;
        198 : data_i <= 16'h04C7;
        199 : data_i <= 16'h04CD;
        200 : data_i <= 16'h04CF;
        201 : data_i <= 16'h04D5;
        202 : data_i <= 16'h04E1;
        203 : data_i <= 16'h04EB;
        204 : data_i <= 16'h04FD;
        205 : data_i <= 16'h04FF;
        206 : data_i <= 16'h0503;
        207 : data_i <= 16'h0509;
        208 : data_i <= 16'h050B;
        209 : data_i <= 16'h0511;
        210 : data_i <= 16'h0515;
        211 : data_i <= 16'h0517;
        212 : data_i <= 16'h051B;
        213 : data_i <= 16'h0527;
        214 : data_i <= 16'h0529;
        215 : data_i <= 16'h052F;
        216 : data_i <= 16'h0551;
        217 : data_i <= 16'h0557;
        218 : data_i <= 16'h055D;
        219 : data_i <= 16'h0565;
        220 : data_i <= 16'h0577;
        221 : data_i <= 16'h0581;
        222 : data_i <= 16'h058F;
        223 : data_i <= 16'h0593;
        224 : data_i <= 16'h0595;
        225 : data_i <= 16'h0599;
        226 : data_i <= 16'h059F;
        227 : data_i <= 16'h05A7;
        228 : data_i <= 16'h05AB;
        229 : data_i <= 16'h05AD;
        230 : data_i <= 16'h05B3;
        231 : data_i <= 16'h05BF;
        232 : data_i <= 16'h05C9;
        233 : data_i <= 16'h05CB;
        234 : data_i <= 16'h05CF;
        235 : data_i <= 16'h05D1;
        236 : data_i <= 16'h05D5;
        237 : data_i <= 16'h05DB;
        238 : data_i <= 16'h05E7;
        239 : data_i <= 16'h05F3;
        240 : data_i <= 16'h05FB;
        241 : data_i <= 16'h0607;
        242 : data_i <= 16'h060D;
        243 : data_i <= 16'h0611;
        244 : data_i <= 16'h0617;
        245 : data_i <= 16'h061F;
        246 : data_i <= 16'h0623;
        247 : data_i <= 16'h062B;
        248 : data_i <= 16'h062F;
        249 : data_i <= 16'h063D;
        250 : data_i <= 16'h0641;
        251 : data_i <= 16'h0647;
        252 : data_i <= 16'h0649;
        253 : data_i <= 16'h064D;
        254 : data_i <= 16'h0653;
        255 : data_i <= 16'h0655;
        256 : data_i <= 16'h065B;
        257 : data_i <= 16'h0665;
        258 : data_i <= 16'h0679;
        259 : data_i <= 16'h067F;
        260 : data_i <= 16'h0683;
        261 : data_i <= 16'h0685;
        262 : data_i <= 16'h069D;
        263 : data_i <= 16'h06A1;
        264 : data_i <= 16'h06A3;
        265 : data_i <= 16'h06AD;
        266 : data_i <= 16'h06B9;
        267 : data_i <= 16'h06BB;
        268 : data_i <= 16'h06C5;
        269 : data_i <= 16'h06CD;
        270 : data_i <= 16'h06D3;
        271 : data_i <= 16'h06D9;
        272 : data_i <= 16'h06DF;
        273 : data_i <= 16'h06F1;
        274 : data_i <= 16'h06F7;
        275 : data_i <= 16'h06FB;
        276 : data_i <= 16'h06FD;
        277 : data_i <= 16'h0709;
        278 : data_i <= 16'h0713;
        279 : data_i <= 16'h071F;
        280 : data_i <= 16'h0727;
        281 : data_i <= 16'h0737;
        282 : data_i <= 16'h0745;
        283 : data_i <= 16'h074B;
        284 : data_i <= 16'h074F;
        285 : data_i <= 16'h0751;
        286 : data_i <= 16'h0755;
        287 : data_i <= 16'h0757;
        288 : data_i <= 16'h0761;
        289 : data_i <= 16'h076D;
        290 : data_i <= 16'h0773;
        291 : data_i <= 16'h0779;
        292 : data_i <= 16'h078B;
        293 : data_i <= 16'h078D;
        294 : data_i <= 16'h079D;
        295 : data_i <= 16'h079F;
        296 : data_i <= 16'h07B5;
        297 : data_i <= 16'h07BB;
        298 : data_i <= 16'h07C3;
        299 : data_i <= 16'h07C9;
        300 : data_i <= 16'h07CD;
        301 : data_i <= 16'h07CF;
        302 : data_i <= 16'h07D3;
        303 : data_i <= 16'h07DB;
        304 : data_i <= 16'h07E1;
        305 : data_i <= 16'h07EB;
        306 : data_i <= 16'h07ED;
        307 : data_i <= 16'h07F7;
        308 : data_i <= 16'h0805;
        309 : data_i <= 16'h080F;
        310 : data_i <= 16'h0815;
        311 : data_i <= 16'h0821;
        312 : data_i <= 16'h0823;
        313 : data_i <= 16'h0827;
        314 : data_i <= 16'h0829;
        315 : data_i <= 16'h0833;
        316 : data_i <= 16'h083F;
        317 : data_i <= 16'h0841;
        318 : data_i <= 16'h0851;
        319 : data_i <= 16'h0853;
        320 : data_i <= 16'h0859;
        321 : data_i <= 16'h085D;
        322 : data_i <= 16'h085F;
        323 : data_i <= 16'h0869;
        324 : data_i <= 16'h0871;
        325 : data_i <= 16'h0883;
        326 : data_i <= 16'h089B;
        327 : data_i <= 16'h089F;
        328 : data_i <= 16'h08A5;
        329 : data_i <= 16'h08AD;
        330 : data_i <= 16'h08BD;
        331 : data_i <= 16'h08BF;
        332 : data_i <= 16'h08C3;
        333 : data_i <= 16'h08CB;
        334 : data_i <= 16'h08DB;
        335 : data_i <= 16'h08DD;
        336 : data_i <= 16'h08E1;
        337 : data_i <= 16'h08E9;
        338 : data_i <= 16'h08EF;
        339 : data_i <= 16'h08F5;
        340 : data_i <= 16'h08F9;
        341 : data_i <= 16'h0905;
        342 : data_i <= 16'h0907;
        343 : data_i <= 16'h091D;
        344 : data_i <= 16'h0923;
        345 : data_i <= 16'h0925;
        346 : data_i <= 16'h092B;
        347 : data_i <= 16'h092F;
        348 : data_i <= 16'h0935;
        349 : data_i <= 16'h0943;
        350 : data_i <= 16'h0949;
        351 : data_i <= 16'h094D;
        352 : data_i <= 16'h094F;
        353 : data_i <= 16'h0955;
        354 : data_i <= 16'h0959;
        355 : data_i <= 16'h095F;
        356 : data_i <= 16'h096B;
        357 : data_i <= 16'h0971;
        358 : data_i <= 16'h0977;
        359 : data_i <= 16'h0985;
        360 : data_i <= 16'h0989;
        361 : data_i <= 16'h098F;
        362 : data_i <= 16'h099B;
        363 : data_i <= 16'h09A3;
        364 : data_i <= 16'h09A9;
        365 : data_i <= 16'h09AD;
        366 : data_i <= 16'h09C7;
        367 : data_i <= 16'h09D9;
        368 : data_i <= 16'h09E3;
        369 : data_i <= 16'h09EB;
        370 : data_i <= 16'h09EF;
        371 : data_i <= 16'h09F5;
        372 : data_i <= 16'h09F7;
        373 : data_i <= 16'h09FD;
        374 : data_i <= 16'h0A13;
        375 : data_i <= 16'h0A1F;
        376 : data_i <= 16'h0A21;
        377 : data_i <= 16'h0A31;
        378 : data_i <= 16'h0A39;
        379 : data_i <= 16'h0A3D;
        380 : data_i <= 16'h0A49;
        381 : data_i <= 16'h0A57;
        382 : data_i <= 16'h0A61;
        383 : data_i <= 16'h0A63;
        384 : data_i <= 16'h0A67;
        385 : data_i <= 16'h0A6F;
        386 : data_i <= 16'h0A75;
        387 : data_i <= 16'h0A7B;
        388 : data_i <= 16'h0A7F;
        389 : data_i <= 16'h0A81;
        390 : data_i <= 16'h0A85;
        391 : data_i <= 16'h0A8B;
        392 : data_i <= 16'h0A93;
        393 : data_i <= 16'h0A97;
        394 : data_i <= 16'h0A99;
        395 : data_i <= 16'h0A9F;
        396 : data_i <= 16'h0AA9;
        397 : data_i <= 16'h0AAB;
        398 : data_i <= 16'h0AB5;
        399 : data_i <= 16'h0ABD;
        400 : data_i <= 16'h0AC1;
        401 : data_i <= 16'h0ACF;
        402 : data_i <= 16'h0AD9;
        403 : data_i <= 16'h0AE5;
        404 : data_i <= 16'h0AE7;
        405 : data_i <= 16'h0AED;
        406 : data_i <= 16'h0AF1;
        407 : data_i <= 16'h0AF3;
        408 : data_i <= 16'h0B03;
        409 : data_i <= 16'h0B11;
        410 : data_i <= 16'h0B15;
        411 : data_i <= 16'h0B1B;
        412 : data_i <= 16'h0B23;
        413 : data_i <= 16'h0B29;
        414 : data_i <= 16'h0B2D;
        415 : data_i <= 16'h0B3F;
        416 : data_i <= 16'h0B47;
        417 : data_i <= 16'h0B51;
        418 : data_i <= 16'h0B57;
        419 : data_i <= 16'h0B5D;
        420 : data_i <= 16'h0B65;
        421 : data_i <= 16'h0B6F;
        422 : data_i <= 16'h0B7B;
        423 : data_i <= 16'h0B89;
        424 : data_i <= 16'h0B8D;
        425 : data_i <= 16'h0B93;
        426 : data_i <= 16'h0B99;
        427 : data_i <= 16'h0B9B;
        428 : data_i <= 16'h0BB7;
        429 : data_i <= 16'h0BB9;
        430 : data_i <= 16'h0BC3;
        431 : data_i <= 16'h0BCB;
        432 : data_i <= 16'h0BCF;
        433 : data_i <= 16'h0BDD;
        434 : data_i <= 16'h0BE1;
        435 : data_i <= 16'h0BE9;
        436 : data_i <= 16'h0BF5;
        437 : data_i <= 16'h0BFB;
        438 : data_i <= 16'h0C07;
        439 : data_i <= 16'h0C0B;
        440 : data_i <= 16'h0C11;
        441 : data_i <= 16'h0C25;
        442 : data_i <= 16'h0C2F;
        443 : data_i <= 16'h0C31;
        444 : data_i <= 16'h0C41;
        445 : data_i <= 16'h0C5B;
        446 : data_i <= 16'h0C5F;
        447 : data_i <= 16'h0C61;
        448 : data_i <= 16'h0C6D;
        449 : data_i <= 16'h0C73;
        450 : data_i <= 16'h0C77;
        451 : data_i <= 16'h0C83;
        452 : data_i <= 16'h0C89;
        453 : data_i <= 16'h0C91;
        454 : data_i <= 16'h0C95;
        455 : data_i <= 16'h0C9D;
        456 : data_i <= 16'h0CB3;
        457 : data_i <= 16'h0CB5;
        458 : data_i <= 16'h0CB9;
        459 : data_i <= 16'h0CBB;
        460 : data_i <= 16'h0CC7;
        461 : data_i <= 16'h0CE3;
        462 : data_i <= 16'h0CE5;
        463 : data_i <= 16'h0CEB;
        464 : data_i <= 16'h0CF1;
        465 : data_i <= 16'h0CF7;
        466 : data_i <= 16'h0CFB;
        467 : data_i <= 16'h0D01;
        468 : data_i <= 16'h0D03;
        469 : data_i <= 16'h0D0F;
        470 : data_i <= 16'h0D13;
        471 : data_i <= 16'h0D1F;
        472 : data_i <= 16'h0D21;
        473 : data_i <= 16'h0D2B;
        474 : data_i <= 16'h0D2D;
        475 : data_i <= 16'h0D3D;
        476 : data_i <= 16'h0D3F;
        477 : data_i <= 16'h0D4F;
        478 : data_i <= 16'h0D55;
        479 : data_i <= 16'h0D69;
        480 : data_i <= 16'h0D79;
        481 : data_i <= 16'h0D81;
        482 : data_i <= 16'h0D85;
        483 : data_i <= 16'h0D87;
        484 : data_i <= 16'h0D8B;
        485 : data_i <= 16'h0D8D;
        486 : data_i <= 16'h0DA3;
        487 : data_i <= 16'h0DAB;
        488 : data_i <= 16'h0DB7;
        489 : data_i <= 16'h0DBD;
        490 : data_i <= 16'h0DC7;
        491 : data_i <= 16'h0DC9;
        492 : data_i <= 16'h0DCD;
        493 : data_i <= 16'h0DD3;
        494 : data_i <= 16'h0DD5;
        495 : data_i <= 16'h0DDB;
        496 : data_i <= 16'h0DE5;
        497 : data_i <= 16'h0DE7;
        498 : data_i <= 16'h0DF3;
        499 : data_i <= 16'h0DFD;
        500 : data_i <= 16'h0DFF;
        501 : data_i <= 16'h0E09;
        502 : data_i <= 16'h0E17;
        503 : data_i <= 16'h0E1D;
        504 : data_i <= 16'h0E21;
        505 : data_i <= 16'h0E27;
        506 : data_i <= 16'h0E2F;
        507 : data_i <= 16'h0E35;
        508 : data_i <= 16'h0E3B;
        509 : data_i <= 16'h0E4B;
        510 : data_i <= 16'h0E57;
        511 : data_i <= 16'h0E59;
        512 : data_i <= 16'h0E5D;
        513 : data_i <= 16'h0E6B;
        514 : data_i <= 16'h0E71;
        515 : data_i <= 16'h0E75;
        516 : data_i <= 16'h0E7D;
        517 : data_i <= 16'h0E87;
        518 : data_i <= 16'h0E8F;
        519 : data_i <= 16'h0E95;
        520 : data_i <= 16'h0E9B;
        521 : data_i <= 16'h0EB1;
        522 : data_i <= 16'h0EB7;
        523 : data_i <= 16'h0EB9;
        524 : data_i <= 16'h0EC3;
        525 : data_i <= 16'h0ED1;
        526 : data_i <= 16'h0ED5;
        527 : data_i <= 16'h0EDB;
        528 : data_i <= 16'h0EED;
        529 : data_i <= 16'h0EEF;
        530 : data_i <= 16'h0EF9;
        531 : data_i <= 16'h0F07;
        532 : data_i <= 16'h0F0B;
        533 : data_i <= 16'h0F0D;
        534 : data_i <= 16'h0F17;
        535 : data_i <= 16'h0F25;
        536 : data_i <= 16'h0F29;
        537 : data_i <= 16'h0F31;
        538 : data_i <= 16'h0F43;
        539 : data_i <= 16'h0F47;
        540 : data_i <= 16'h0F4D;
        541 : data_i <= 16'h0F4F;
        542 : data_i <= 16'h0F53;
        543 : data_i <= 16'h0F59;
        544 : data_i <= 16'h0F5B;
        545 : data_i <= 16'h0F67;
        546 : data_i <= 16'h0F6B;
        547 : data_i <= 16'h0F7F;
        548 : data_i <= 16'h0F95;
        549 : data_i <= 16'h0FA1;
        550 : data_i <= 16'h0FA3;
        551 : data_i <= 16'h0FA7;
        552 : data_i <= 16'h0FAD;
        553 : data_i <= 16'h0FB3;
        554 : data_i <= 16'h0FB5;
        555 : data_i <= 16'h0FBB;
        556 : data_i <= 16'h0FD1;
        557 : data_i <= 16'h0FD3;
        558 : data_i <= 16'h0FD9;
        559 : data_i <= 16'h0FE9;
        560 : data_i <= 16'h0FEF;
        561 : data_i <= 16'h0FFB;
        562 : data_i <= 16'h0FFD;
        563 : data_i <= 16'h1003;
        564 : data_i <= 16'h100F;
        565 : data_i <= 16'h101F;
        566 : data_i <= 16'h1021;
        567 : data_i <= 16'h1025;
        568 : data_i <= 16'h102B;
        569 : data_i <= 16'h1039;
        570 : data_i <= 16'h103D;
        571 : data_i <= 16'h103F;
        572 : data_i <= 16'h1051;
        573 : data_i <= 16'h1069;
        574 : data_i <= 16'h1073;
        575 : data_i <= 16'h1079;
        576 : data_i <= 16'h107B;
        577 : data_i <= 16'h1085;
        578 : data_i <= 16'h1087;
        579 : data_i <= 16'h1091;
        580 : data_i <= 16'h1093;
        581 : data_i <= 16'h109D;
        582 : data_i <= 16'h10A3;
        583 : data_i <= 16'h10A5;
        584 : data_i <= 16'h10AF;
        585 : data_i <= 16'h10B1;
        586 : data_i <= 16'h10BB;
        587 : data_i <= 16'h10C1;
        588 : data_i <= 16'h10C9;
        589 : data_i <= 16'h10E7;
        590 : data_i <= 16'h10F1;
        591 : data_i <= 16'h10F3;
        592 : data_i <= 16'h10FD;
        593 : data_i <= 16'h1105;
        594 : data_i <= 16'h110B;
        595 : data_i <= 16'h1115;
        596 : data_i <= 16'h1127;
        597 : data_i <= 16'h112D;
        598 : data_i <= 16'h1139;
        599 : data_i <= 16'h1145;
        600 : data_i <= 16'h1147;
        601 : data_i <= 16'h1159;
        602 : data_i <= 16'h115F;
        603 : data_i <= 16'h1163;
        604 : data_i <= 16'h1169;
        605 : data_i <= 16'h116F;
        606 : data_i <= 16'h1181;
        607 : data_i <= 16'h1183;
        608 : data_i <= 16'h118D;
        609 : data_i <= 16'h119B;
        610 : data_i <= 16'h11A1;
        611 : data_i <= 16'h11A5;
        612 : data_i <= 16'h11A7;
        613 : data_i <= 16'h11AB;
        614 : data_i <= 16'h11C3;
        615 : data_i <= 16'h11C5;
        616 : data_i <= 16'h11D1;
        617 : data_i <= 16'h11D7;
        618 : data_i <= 16'h11E7;
        619 : data_i <= 16'h11EF;
        620 : data_i <= 16'h11F5;
        621 : data_i <= 16'h11FB;
        622 : data_i <= 16'h120D;
        623 : data_i <= 16'h121D;
        624 : data_i <= 16'h121F;
        625 : data_i <= 16'h1223;
        626 : data_i <= 16'h1229;
        627 : data_i <= 16'h122B;
        628 : data_i <= 16'h1231;
        629 : data_i <= 16'h1237;
        630 : data_i <= 16'h1241;
        631 : data_i <= 16'h1247;
        632 : data_i <= 16'h1253;
        633 : data_i <= 16'h125F;
        634 : data_i <= 16'h1271;
        635 : data_i <= 16'h1273;
        636 : data_i <= 16'h1279;
        637 : data_i <= 16'h127D;
        638 : data_i <= 16'h128F;
        639 : data_i <= 16'h1297;
        640 : data_i <= 16'h12AF;
        641 : data_i <= 16'h12B3;
        642 : data_i <= 16'h12B5;
        643 : data_i <= 16'h12B9;
        644 : data_i <= 16'h12BF;
        645 : data_i <= 16'h12C1;
        646 : data_i <= 16'h12CD;
        647 : data_i <= 16'h12D1;
        648 : data_i <= 16'h12DF;
        649 : data_i <= 16'h12FD;
        650 : data_i <= 16'h1307;
        651 : data_i <= 16'h130D;
        652 : data_i <= 16'h1319;
        653 : data_i <= 16'h1327;
        654 : data_i <= 16'h132D;
        655 : data_i <= 16'h1337;
        656 : data_i <= 16'h1343;
        657 : data_i <= 16'h1345;
        658 : data_i <= 16'h1349;
        659 : data_i <= 16'h134F;
        660 : data_i <= 16'h1357;
        661 : data_i <= 16'h135D;
        662 : data_i <= 16'h1367;
        663 : data_i <= 16'h1369;
        664 : data_i <= 16'h136D;
        665 : data_i <= 16'h137B;
        666 : data_i <= 16'h1381;
        667 : data_i <= 16'h1387;
        668 : data_i <= 16'h138B;
        669 : data_i <= 16'h1391;
        670 : data_i <= 16'h1393;
        671 : data_i <= 16'h139D;
        672 : data_i <= 16'h139F;
        673 : data_i <= 16'h13AF;
        674 : data_i <= 16'h13BB;
        675 : data_i <= 16'h13C3;
        676 : data_i <= 16'h13D5;
        677 : data_i <= 16'h13D9;
        678 : data_i <= 16'h13DF;
        679 : data_i <= 16'h13EB;
        680 : data_i <= 16'h13ED;
        681 : data_i <= 16'h13F3;
        682 : data_i <= 16'h13F9;
        683 : data_i <= 16'h13FF;
        684 : data_i <= 16'h141B;
        685 : data_i <= 16'h1421;
        686 : data_i <= 16'h142F;
        687 : data_i <= 16'h1433;
        688 : data_i <= 16'h143B;
        689 : data_i <= 16'h1445;
        690 : data_i <= 16'h144D;
        691 : data_i <= 16'h1459;
        692 : data_i <= 16'h146B;
        693 : data_i <= 16'h146F;
        694 : data_i <= 16'h1471;
        695 : data_i <= 16'h1475;
        696 : data_i <= 16'h148D;
        697 : data_i <= 16'h1499;
        698 : data_i <= 16'h149F;
        699 : data_i <= 16'h14A1;
        700 : data_i <= 16'h14B1;
        701 : data_i <= 16'h14B7;
        702 : data_i <= 16'h14BD;
        703 : data_i <= 16'h14CB;
        704 : data_i <= 16'h14D5;
        705 : data_i <= 16'h14E3;
        706 : data_i <= 16'h14E7;
        707 : data_i <= 16'h1505;
        708 : data_i <= 16'h150B;
        709 : data_i <= 16'h1511;
        710 : data_i <= 16'h1517;
        711 : data_i <= 16'h151F;
        712 : data_i <= 16'h1525;
        713 : data_i <= 16'h1529;
        714 : data_i <= 16'h152B;
        715 : data_i <= 16'h1537;
        716 : data_i <= 16'h153D;
        717 : data_i <= 16'h1541;
        718 : data_i <= 16'h1543;
        719 : data_i <= 16'h1549;
        720 : data_i <= 16'h155F;
        721 : data_i <= 16'h1565;
        722 : data_i <= 16'h1567;
        723 : data_i <= 16'h156B;
        724 : data_i <= 16'h157D;
        725 : data_i <= 16'h157F;
        726 : data_i <= 16'h1583;
        727 : data_i <= 16'h158F;
        728 : data_i <= 16'h1591;
        729 : data_i <= 16'h1597;
        730 : data_i <= 16'h159B;
        731 : data_i <= 16'h15B5;
        732 : data_i <= 16'h15BB;
        733 : data_i <= 16'h15C1;
        734 : data_i <= 16'h15C5;
        735 : data_i <= 16'h15CD;
        736 : data_i <= 16'h15D7;
        737 : data_i <= 16'h15F7;
        738 : data_i <= 16'h1607;
        739 : data_i <= 16'h1609;
        740 : data_i <= 16'h160F;
        741 : data_i <= 16'h1613;
        742 : data_i <= 16'h1615;
        743 : data_i <= 16'h1619;
        744 : data_i <= 16'h161B;
        745 : data_i <= 16'h1625;
        746 : data_i <= 16'h1633;
        747 : data_i <= 16'h1639;
        748 : data_i <= 16'h163D;
        749 : data_i <= 16'h1645;
        750 : data_i <= 16'h164F;
        751 : data_i <= 16'h1655;
        752 : data_i <= 16'h1669;
        753 : data_i <= 16'h166D;
        754 : data_i <= 16'h166F;
        755 : data_i <= 16'h1675;
        756 : data_i <= 16'h1693;
        757 : data_i <= 16'h1697;
        758 : data_i <= 16'h169F;
        759 : data_i <= 16'h16A9;
        760 : data_i <= 16'h16AF;
        761 : data_i <= 16'h16B5;
        762 : data_i <= 16'h16BD;
        763 : data_i <= 16'h16C3;
        764 : data_i <= 16'h16CF;
        765 : data_i <= 16'h16D3;
        766 : data_i <= 16'h16D9;
        767 : data_i <= 16'h16DB;
        768 : data_i <= 16'h16E1;
        769 : data_i <= 16'h16E5;
        770 : data_i <= 16'h16EB;
        771 : data_i <= 16'h16ED;
        772 : data_i <= 16'h16F7;
        773 : data_i <= 16'h16F9;
        774 : data_i <= 16'h1709;
        775 : data_i <= 16'h170F;
        776 : data_i <= 16'h1723;
        777 : data_i <= 16'h1727;
        778 : data_i <= 16'h1733;
        779 : data_i <= 16'h1741;
        780 : data_i <= 16'h175D;
        781 : data_i <= 16'h1763;
        782 : data_i <= 16'h1777;
        783 : data_i <= 16'h177B;
        784 : data_i <= 16'h178D;
        785 : data_i <= 16'h1795;
        786 : data_i <= 16'h179B;
        787 : data_i <= 16'h179F;
        788 : data_i <= 16'h17A5;
        789 : data_i <= 16'h17B3;
        790 : data_i <= 16'h17B9;
        791 : data_i <= 16'h17BF;
        792 : data_i <= 16'h17C9;
        793 : data_i <= 16'h17CB;
        794 : data_i <= 16'h17D5;
        795 : data_i <= 16'h17E1;
        796 : data_i <= 16'h17E9;
        797 : data_i <= 16'h17F3;
        798 : data_i <= 16'h17F5;
        799 : data_i <= 16'h17FF;
        800 : data_i <= 16'h1807;
        801 : data_i <= 16'h1813;
        802 : data_i <= 16'h181D;
        803 : data_i <= 16'h1835;
        804 : data_i <= 16'h1837;
        805 : data_i <= 16'h183B;
        806 : data_i <= 16'h1843;
        807 : data_i <= 16'h1849;
        808 : data_i <= 16'h184D;
        809 : data_i <= 16'h1855;
        810 : data_i <= 16'h1867;
        811 : data_i <= 16'h1871;
        812 : data_i <= 16'h1877;
        813 : data_i <= 16'h187D;
        814 : data_i <= 16'h187F;
        815 : data_i <= 16'h1885;
        816 : data_i <= 16'h188F;
        817 : data_i <= 16'h189B;
        818 : data_i <= 16'h189D;
        819 : data_i <= 16'h18A7;
        820 : data_i <= 16'h18AD;
        821 : data_i <= 16'h18B3;
        822 : data_i <= 16'h18B9;
        823 : data_i <= 16'h18C1;
        824 : data_i <= 16'h18C7;
        825 : data_i <= 16'h18D1;
        826 : data_i <= 16'h18D7;
        827 : data_i <= 16'h18D9;
        828 : data_i <= 16'h18DF;
        829 : data_i <= 16'h18E5;
        830 : data_i <= 16'h18EB;
        831 : data_i <= 16'h18F5;
        832 : data_i <= 16'h18FD;
        833 : data_i <= 16'h1915;
        834 : data_i <= 16'h191B;
        835 : data_i <= 16'h1931;
        836 : data_i <= 16'h1933;
        837 : data_i <= 16'h1945;
        838 : data_i <= 16'h1949;
        839 : data_i <= 16'h1951;
        840 : data_i <= 16'h195B;
        841 : data_i <= 16'h1979;
        842 : data_i <= 16'h1981;
        843 : data_i <= 16'h1993;
        844 : data_i <= 16'h1997;
        845 : data_i <= 16'h1999;
        846 : data_i <= 16'h19A3;
        847 : data_i <= 16'h19A9;
        848 : data_i <= 16'h19AB;
        849 : data_i <= 16'h19B1;
        850 : data_i <= 16'h19B5;
        851 : data_i <= 16'h19C7;
        852 : data_i <= 16'h19CF;
        853 : data_i <= 16'h19DB;
        854 : data_i <= 16'h19ED;
        855 : data_i <= 16'h19FD;
        856 : data_i <= 16'h1A03;
        857 : data_i <= 16'h1A05;
        858 : data_i <= 16'h1A11;
        859 : data_i <= 16'h1A17;
        860 : data_i <= 16'h1A21;
        861 : data_i <= 16'h1A23;
        862 : data_i <= 16'h1A2D;
        863 : data_i <= 16'h1A2F;
        864 : data_i <= 16'h1A35;
        865 : data_i <= 16'h1A3F;
        866 : data_i <= 16'h1A4D;
        867 : data_i <= 16'h1A51;
        868 : data_i <= 16'h1A69;
        869 : data_i <= 16'h1A6B;
        870 : data_i <= 16'h1A7B;
        871 : data_i <= 16'h1A7D;
        872 : data_i <= 16'h1A87;
        873 : data_i <= 16'h1A89;
        874 : data_i <= 16'h1A93;
        875 : data_i <= 16'h1AA7;
        876 : data_i <= 16'h1AAB;
        877 : data_i <= 16'h1AAD;
        878 : data_i <= 16'h1AB1;
        879 : data_i <= 16'h1AB9;
        880 : data_i <= 16'h1AC9;
        881 : data_i <= 16'h1ACF;
        882 : data_i <= 16'h1AD5;
        883 : data_i <= 16'h1AD7;
        884 : data_i <= 16'h1AE3;
        885 : data_i <= 16'h1AF3;
        886 : data_i <= 16'h1AFB;
        887 : data_i <= 16'h1AFF;
        888 : data_i <= 16'h1B05;
        889 : data_i <= 16'h1B23;
        890 : data_i <= 16'h1B25;
        891 : data_i <= 16'h1B2F;
        892 : data_i <= 16'h1B31;
        893 : data_i <= 16'h1B37;
        894 : data_i <= 16'h1B3B;
        895 : data_i <= 16'h1B41;
        896 : data_i <= 16'h1B47;
        897 : data_i <= 16'h1B4F;
        898 : data_i <= 16'h1B55;
        899 : data_i <= 16'h1B59;
        900 : data_i <= 16'h1B65;
        901 : data_i <= 16'h1B6B;
        902 : data_i <= 16'h1B73;
        903 : data_i <= 16'h1B7F;
        904 : data_i <= 16'h1B83;
        905 : data_i <= 16'h1B91;
        906 : data_i <= 16'h1B9D;
        907 : data_i <= 16'h1BA7;
        908 : data_i <= 16'h1BBF;
        909 : data_i <= 16'h1BC5;
        910 : data_i <= 16'h1BD1;
        911 : data_i <= 16'h1BD7;
        912 : data_i <= 16'h1BD9;
        913 : data_i <= 16'h1BEF;
        914 : data_i <= 16'h1BF7;
        915 : data_i <= 16'h1C09;
        916 : data_i <= 16'h1C13;
        917 : data_i <= 16'h1C19;
        918 : data_i <= 16'h1C27;
        919 : data_i <= 16'h1C2B;
        920 : data_i <= 16'h1C2D;
        921 : data_i <= 16'h1C33;
        922 : data_i <= 16'h1C3D;
        923 : data_i <= 16'h1C45;
        924 : data_i <= 16'h1C4B;
        925 : data_i <= 16'h1C4F;
        926 : data_i <= 16'h1C55;
        927 : data_i <= 16'h1C73;
        928 : data_i <= 16'h1C81;
        929 : data_i <= 16'h1C8B;
        930 : data_i <= 16'h1C8D;
        931 : data_i <= 16'h1C99;
        932 : data_i <= 16'h1CA3;
        933 : data_i <= 16'h1CA5;
        934 : data_i <= 16'h1CB5;
        935 : data_i <= 16'h1CB7;
        936 : data_i <= 16'h1CC9;
        937 : data_i <= 16'h1CE1;
        938 : data_i <= 16'h1CF3;
        939 : data_i <= 16'h1CF9;
        940 : data_i <= 16'h1D09;
        941 : data_i <= 16'h1D1B;
        942 : data_i <= 16'h1D21;
        943 : data_i <= 16'h1D23;
        944 : data_i <= 16'h1D35;
        945 : data_i <= 16'h1D39;
        946 : data_i <= 16'h1D3F;
        947 : data_i <= 16'h1D41;
        948 : data_i <= 16'h1D4B;
        949 : data_i <= 16'h1D53;
        950 : data_i <= 16'h1D5D;
        951 : data_i <= 16'h1D63;
        952 : data_i <= 16'h1D69;
        953 : data_i <= 16'h1D71;
        954 : data_i <= 16'h1D75;
        955 : data_i <= 16'h1D7B;
        956 : data_i <= 16'h1D7D;
        957 : data_i <= 16'h1D87;
        958 : data_i <= 16'h1D89;
        959 : data_i <= 16'h1D95;
        960 : data_i <= 16'h1D99;
        961 : data_i <= 16'h1D9F;
        962 : data_i <= 16'h1DA5;
        963 : data_i <= 16'h1DA7;
        964 : data_i <= 16'h1DB3;
        965 : data_i <= 16'h1DB7;
        966 : data_i <= 16'h1DC5;
        967 : data_i <= 16'h1DD7;
        968 : data_i <= 16'h1DDB;
        969 : data_i <= 16'h1DE1;
        970 : data_i <= 16'h1DF5;
        971 : data_i <= 16'h1DF9;
        972 : data_i <= 16'h1E01;
        973 : data_i <= 16'h1E07;
        974 : data_i <= 16'h1E0B;
        975 : data_i <= 16'h1E13;
        976 : data_i <= 16'h1E17;
        977 : data_i <= 16'h1E25;
        978 : data_i <= 16'h1E2B;
        979 : data_i <= 16'h1E2F;
        980 : data_i <= 16'h1E3D;
        981 : data_i <= 16'h1E49;
        982 : data_i <= 16'h1E4D;
        983 : data_i <= 16'h1E4F;
        984 : data_i <= 16'h1E6D;
        985 : data_i <= 16'h1E71;
        986 : data_i <= 16'h1E89;
        987 : data_i <= 16'h1E8F;
        988 : data_i <= 16'h1E95;
        989 : data_i <= 16'h1EA1;
        990 : data_i <= 16'h1EAD;
        991 : data_i <= 16'h1EBB;
        992 : data_i <= 16'h1EC1;
        993 : data_i <= 16'h1EC5;
        994 : data_i <= 16'h1EC7;
        995 : data_i <= 16'h1ECB;
        996 : data_i <= 16'h1EDD;
        997 : data_i <= 16'h1EE3;
        998 : data_i <= 16'h1EEF;
        999 : data_i <= 16'h1EF7;
        1000 : data_i <= 16'h1EFD;
        1001 : data_i <= 16'h1F01;
        1002 : data_i <= 16'h1F0D;
        1003 : data_i <= 16'h1F0F;
        1004 : data_i <= 16'h1F1B;
        1005 : data_i <= 16'h1F39;
        1006 : data_i <= 16'h1F49;
        1007 : data_i <= 16'h1F4B;
        1008 : data_i <= 16'h1F51;
        1009 : data_i <= 16'h1F67;
        1010 : data_i <= 16'h1F75;
        1011 : data_i <= 16'h1F7B;
        1012 : data_i <= 16'h1F85;
        1013 : data_i <= 16'h1F91;
        1014 : data_i <= 16'h1F97;
        1015 : data_i <= 16'h1F99;
        1016 : data_i <= 16'h1F9D;
        1017 : data_i <= 16'h1FA5;
        1018 : data_i <= 16'h1FAF;
        1019 : data_i <= 16'h1FB5;
        1020 : data_i <= 16'h1FBB;
        1021 : data_i <= 16'h1FD3;
        1022 : data_i <= 16'h1FE1;
        1023 : data_i <= 16'h1FE7;
        1024 : data_i <= 16'h1FEB;
        1025 : data_i <= 16'h1FF3;
        1026 : data_i <= 16'h1FFF;
        1027 : data_i <= 16'h2011;
        1028 : data_i <= 16'h201B;
        1029 : data_i <= 16'h201D;
        1030 : data_i <= 16'h2027;
        1031 : data_i <= 16'h2029;
        1032 : data_i <= 16'h202D;
        1033 : data_i <= 16'h2033;
        1034 : data_i <= 16'h2047;
        1035 : data_i <= 16'h204D;
        1036 : data_i <= 16'h2051;
        1037 : data_i <= 16'h205F;
        1038 : data_i <= 16'h2063;
        1039 : data_i <= 16'h2065;
        1040 : data_i <= 16'h2069;
        1041 : data_i <= 16'h2077;
        1042 : data_i <= 16'h207D;
        1043 : data_i <= 16'h2089;
        1044 : data_i <= 16'h20A1;
        1045 : data_i <= 16'h20AB;
        1046 : data_i <= 16'h20B1;
        1047 : data_i <= 16'h20B9;
        1048 : data_i <= 16'h20C3;
        1049 : data_i <= 16'h20C5;
        1050 : data_i <= 16'h20E3;
        1051 : data_i <= 16'h20E7;
        1052 : data_i <= 16'h20ED;
        1053 : data_i <= 16'h20EF;
        1054 : data_i <= 16'h20FB;
        1055 : data_i <= 16'h20FF;
        1056 : data_i <= 16'h210D;
        1057 : data_i <= 16'h2113;
        1058 : data_i <= 16'h2135;
        1059 : data_i <= 16'h2141;
        1060 : data_i <= 16'h2149;
        1061 : data_i <= 16'h214F;
        1062 : data_i <= 16'h2159;
        1063 : data_i <= 16'h215B;
        1064 : data_i <= 16'h215F;
        1065 : data_i <= 16'h2173;
        1066 : data_i <= 16'h217D;
        1067 : data_i <= 16'h2185;
        1068 : data_i <= 16'h2195;
        1069 : data_i <= 16'h2197;
        1070 : data_i <= 16'h21A1;
        1071 : data_i <= 16'h21AF;
        1072 : data_i <= 16'h21B3;
        1073 : data_i <= 16'h21B5;
        1074 : data_i <= 16'h21C1;
        1075 : data_i <= 16'h21C7;
        1076 : data_i <= 16'h21D7;
        1077 : data_i <= 16'h21DD;
        1078 : data_i <= 16'h21E5;
        1079 : data_i <= 16'h21E9;
        1080 : data_i <= 16'h21F1;
        1081 : data_i <= 16'h21F5;
        1082 : data_i <= 16'h21FB;
        1083 : data_i <= 16'h2203;
        1084 : data_i <= 16'h2209;
        1085 : data_i <= 16'h220F;
        1086 : data_i <= 16'h221B;
        1087 : data_i <= 16'h2221;
        1088 : data_i <= 16'h2225;
        1089 : data_i <= 16'h222B;
        1090 : data_i <= 16'h2231;
        1091 : data_i <= 16'h2239;
        1092 : data_i <= 16'h224B;
        1093 : data_i <= 16'h224F;
        1094 : data_i <= 16'h2263;
        1095 : data_i <= 16'h2267;
        1096 : data_i <= 16'h2273;
        1097 : data_i <= 16'h2275;
        1098 : data_i <= 16'h227F;
        1099 : data_i <= 16'h2285;
        1100 : data_i <= 16'h2287;
        1101 : data_i <= 16'h2291;
        1102 : data_i <= 16'h229D;
        1103 : data_i <= 16'h229F;
        1104 : data_i <= 16'h22A3;
        1105 : data_i <= 16'h22B7;
        1106 : data_i <= 16'h22BD;
        1107 : data_i <= 16'h22DB;
        1108 : data_i <= 16'h22E1;
        1109 : data_i <= 16'h22E5;
        1110 : data_i <= 16'h22ED;
        1111 : data_i <= 16'h22F7;
        1112 : data_i <= 16'h2303;
        1113 : data_i <= 16'h2309;
        1114 : data_i <= 16'h230B;
        1115 : data_i <= 16'h2327;
        1116 : data_i <= 16'h2329;
        1117 : data_i <= 16'h232F;
        1118 : data_i <= 16'h2333;
        1119 : data_i <= 16'h2335;
        1120 : data_i <= 16'h2345;
        1121 : data_i <= 16'h2351;
        1122 : data_i <= 16'h2353;
        1123 : data_i <= 16'h2359;
        1124 : data_i <= 16'h2363;
        1125 : data_i <= 16'h236B;
        1126 : data_i <= 16'h2383;
        1127 : data_i <= 16'h238F;
        1128 : data_i <= 16'h2395;
        1129 : data_i <= 16'h23A7;
        1130 : data_i <= 16'h23AD;
        1131 : data_i <= 16'h23B1;
        1132 : data_i <= 16'h23BF;
        1133 : data_i <= 16'h23C5;
        1134 : data_i <= 16'h23C9;
        1135 : data_i <= 16'h23D5;
        1136 : data_i <= 16'h23DD;
        1137 : data_i <= 16'h23E3;
        1138 : data_i <= 16'h23EF;
        1139 : data_i <= 16'h23F3;
        1140 : data_i <= 16'h23F9;
        1141 : data_i <= 16'h2405;
        1142 : data_i <= 16'h240B;
        1143 : data_i <= 16'h2417;
        1144 : data_i <= 16'h2419;
        1145 : data_i <= 16'h2429;
        1146 : data_i <= 16'h243D;
        1147 : data_i <= 16'h2441;
        1148 : data_i <= 16'h2443;
        1149 : data_i <= 16'h244D;
        1150 : data_i <= 16'h245F;
        1151 : data_i <= 16'h2467;
        1152 : data_i <= 16'h246B;
        1153 : data_i <= 16'h2479;
        1154 : data_i <= 16'h247D;
        1155 : data_i <= 16'h247F;
        1156 : data_i <= 16'h2485;
        1157 : data_i <= 16'h249B;
        1158 : data_i <= 16'h24A1;
        1159 : data_i <= 16'h24AF;
        1160 : data_i <= 16'h24B5;
        1161 : data_i <= 16'h24BB;
        1162 : data_i <= 16'h24C5;
        1163 : data_i <= 16'h24CB;
        1164 : data_i <= 16'h24CD;
        1165 : data_i <= 16'h24D7;
        1166 : data_i <= 16'h24D9;
        1167 : data_i <= 16'h24DD;
        1168 : data_i <= 16'h24DF;
        1169 : data_i <= 16'h24F5;
        1170 : data_i <= 16'h24F7;
        1171 : data_i <= 16'h24FB;
        1172 : data_i <= 16'h2501;
        1173 : data_i <= 16'h2507;
        1174 : data_i <= 16'h2513;
        1175 : data_i <= 16'h2519;
        1176 : data_i <= 16'h2527;
        1177 : data_i <= 16'h2531;
        1178 : data_i <= 16'h253D;
        1179 : data_i <= 16'h2543;
        1180 : data_i <= 16'h254B;
        1181 : data_i <= 16'h254F;
        1182 : data_i <= 16'h2573;
        1183 : data_i <= 16'h2581;
        1184 : data_i <= 16'h258D;
        1185 : data_i <= 16'h2593;
        1186 : data_i <= 16'h2597;
        1187 : data_i <= 16'h259D;
        1188 : data_i <= 16'h259F;
        1189 : data_i <= 16'h25AB;
        1190 : data_i <= 16'h25B1;
        1191 : data_i <= 16'h25BD;
        1192 : data_i <= 16'h25CD;
        1193 : data_i <= 16'h25CF;
        1194 : data_i <= 16'h25D9;
        1195 : data_i <= 16'h25E1;
        1196 : data_i <= 16'h25F7;
        1197 : data_i <= 16'h25F9;
        1198 : data_i <= 16'h2605;
        1199 : data_i <= 16'h260B;
        1200 : data_i <= 16'h260F;
        1201 : data_i <= 16'h2615;
        1202 : data_i <= 16'h2627;
        1203 : data_i <= 16'h2629;
        1204 : data_i <= 16'h2635;
        1205 : data_i <= 16'h263B;
        1206 : data_i <= 16'h263F;
        1207 : data_i <= 16'h264B;
        1208 : data_i <= 16'h2653;
        1209 : data_i <= 16'h2659;
        1210 : data_i <= 16'h2665;
        1211 : data_i <= 16'h2669;
        1212 : data_i <= 16'h266F;
        1213 : data_i <= 16'h267B;
        1214 : data_i <= 16'h2681;
        1215 : data_i <= 16'h2683;
        1216 : data_i <= 16'h268F;
        1217 : data_i <= 16'h269B;
        1218 : data_i <= 16'h269F;
        1219 : data_i <= 16'h26AD;
        1220 : data_i <= 16'h26B3;
        1221 : data_i <= 16'h26C3;
        1222 : data_i <= 16'h26C9;
        1223 : data_i <= 16'h26CB;
        1224 : data_i <= 16'h26D5;
        1225 : data_i <= 16'h26DD;
        1226 : data_i <= 16'h26EF;
        1227 : data_i <= 16'h26F5;
    endcase
end

assign DATA = data_i;


endmodule    //PRIME_ROM