-- =====================================================================
--  Title       : Prime number ROM
--
--  File Name	: PRIME_ROM.vhd
--  Project     :
--  Block       :
--  Tree        :
--  Designer    : toms74209200 <https://github.com/toms74209200>
--  Created     : 2019/09/22
--  Copyright   : 2019 toms74209200
--  License     : MIT License.
--                http://opensource.org/licenses/mit-license.php
-- =====================================================================
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity PRIME_ROM is
    port(
    -- System --
        CLK     : in    std_logic;                          --(p) Clock

    -- ROM interface --
        ADDRESS : in    std_logic_vector(10 downto 0);      --(p) Address
        DATA    : out   std_logic_vector(15 downto 0)       --(p) Data
        );
end PRIME_ROM;

architecture RTL of PRIME_ROM is

-- Internal signals --
signal data_i           : std_logic_vector(DATA'range);     -- Data

begin
-- ***********************************************************
--  ROM output
-- ***********************************************************
process (CLK) begin
    if (CLK'event and CLK = '1') then
        case (CONV_INTEGER(ADDRESS)) is
            when 0   => data_i <= X"0003";
            when 1   => data_i <= X"0005";
            when 2   => data_i <= X"0007";
            when 3   => data_i <= X"000B";
            when 4   => data_i <= X"000D";
            when 5   => data_i <= X"0011";
            when 6   => data_i <= X"0013";
            when 7   => data_i <= X"0017";
            when 8   => data_i <= X"001D";
            when 9   => data_i <= X"001F";
            when 10  => data_i <= X"0025";
            when 11  => data_i <= X"0029";
            when 12  => data_i <= X"002B";
            when 13  => data_i <= X"002F";
            when 14  => data_i <= X"0035";
            when 15  => data_i <= X"003B";
            when 16  => data_i <= X"003D";
            when 17  => data_i <= X"0043";
            when 18  => data_i <= X"0047";
            when 19  => data_i <= X"0049";
            when 20  => data_i <= X"004F";
            when 21  => data_i <= X"0053";
            when 22  => data_i <= X"0059";
            when 23  => data_i <= X"0061";
            when 24  => data_i <= X"0065";
            when 25  => data_i <= X"0067";
            when 26  => data_i <= X"006B";
            when 27  => data_i <= X"006D";
            when 28  => data_i <= X"0071";
            when 29  => data_i <= X"007F";
            when 30  => data_i <= X"0083";
            when 31  => data_i <= X"0089";
            when 32  => data_i <= X"008B";
            when 33  => data_i <= X"0095";
            when 34  => data_i <= X"0097";
            when 35  => data_i <= X"009D";
            when 36  => data_i <= X"00A3";
            when 37  => data_i <= X"00A7";
            when 38  => data_i <= X"00AD";
            when 39  => data_i <= X"00B3";
            when 40  => data_i <= X"00B5";
            when 41  => data_i <= X"00BF";
            when 42  => data_i <= X"00C1";
            when 43  => data_i <= X"00C5";
            when 44  => data_i <= X"00C7";
            when 45  => data_i <= X"00D3";
            when 46  => data_i <= X"00DF";
            when 47  => data_i <= X"00E3";
            when 48  => data_i <= X"00E5";
            when 49  => data_i <= X"00E9";
            when 50  => data_i <= X"00EF";
            when 51  => data_i <= X"00F1";
            when 52  => data_i <= X"00FB";
            when 53  => data_i <= X"0101";
            when 54  => data_i <= X"0107";
            when 55  => data_i <= X"010D";
            when 56  => data_i <= X"010F";
            when 57  => data_i <= X"0115";
            when 58  => data_i <= X"0119";
            when 59  => data_i <= X"011B";
            when 60  => data_i <= X"0125";
            when 61  => data_i <= X"0133";
            when 62  => data_i <= X"0137";
            when 63  => data_i <= X"0139";
            when 64  => data_i <= X"013D";
            when 65  => data_i <= X"014B";
            when 66  => data_i <= X"0151";
            when 67  => data_i <= X"015B";
            when 68  => data_i <= X"015D";
            when 69  => data_i <= X"0161";
            when 70  => data_i <= X"0167";
            when 71  => data_i <= X"016F";
            when 72  => data_i <= X"0175";
            when 73  => data_i <= X"017B";
            when 74  => data_i <= X"017F";
            when 75  => data_i <= X"0185";
            when 76  => data_i <= X"018D";
            when 77  => data_i <= X"0191";
            when 78  => data_i <= X"0199";
            when 79  => data_i <= X"01A3";
            when 80  => data_i <= X"01A5";
            when 81  => data_i <= X"01AF";
            when 82  => data_i <= X"01B1";
            when 83  => data_i <= X"01B7";
            when 84  => data_i <= X"01BB";
            when 85  => data_i <= X"01C1";
            when 86  => data_i <= X"01C9";
            when 87  => data_i <= X"01CD";
            when 88  => data_i <= X"01CF";
            when 89  => data_i <= X"01D3";
            when 90  => data_i <= X"01DF";
            when 91  => data_i <= X"01E7";
            when 92  => data_i <= X"01EB";
            when 93  => data_i <= X"01F3";
            when 94  => data_i <= X"01F7";
            when 95  => data_i <= X"01FD";
            when 96  => data_i <= X"0209";
            when 97  => data_i <= X"020B";
            when 98  => data_i <= X"021D";
            when 99  => data_i <= X"0223";
            when 100 => data_i <= X"022D";
            when 101 => data_i <= X"0233";
            when 102 => data_i <= X"0239";
            when 103 => data_i <= X"023B";
            when 104 => data_i <= X"0241";
            when 105 => data_i <= X"024B";
            when 106 => data_i <= X"0251";
            when 107 => data_i <= X"0257";
            when 108 => data_i <= X"0259";
            when 109 => data_i <= X"025F";
            when 110 => data_i <= X"0265";
            when 111 => data_i <= X"0269";
            when 112 => data_i <= X"026B";
            when 113 => data_i <= X"0277";
            when 114 => data_i <= X"0281";
            when 115 => data_i <= X"0283";
            when 116 => data_i <= X"0287";
            when 117 => data_i <= X"028D";
            when 118 => data_i <= X"0293";
            when 119 => data_i <= X"0295";
            when 120 => data_i <= X"02A1";
            when 121 => data_i <= X"02A5";
            when 122 => data_i <= X"02AB";
            when 123 => data_i <= X"02B3";
            when 124 => data_i <= X"02BD";
            when 125 => data_i <= X"02C5";
            when 126 => data_i <= X"02CF";
            when 127 => data_i <= X"02D7";
            when 128 => data_i <= X"02DD";
            when 129 => data_i <= X"02E3";
            when 130 => data_i <= X"02E7";
            when 131 => data_i <= X"02EF";
            when 132 => data_i <= X"02F5";
            when 133 => data_i <= X"02F9";
            when 134 => data_i <= X"0301";
            when 135 => data_i <= X"0305";
            when 136 => data_i <= X"0313";
            when 137 => data_i <= X"031D";
            when 138 => data_i <= X"0329";
            when 139 => data_i <= X"032B";
            when 140 => data_i <= X"0335";
            when 141 => data_i <= X"0337";
            when 142 => data_i <= X"033B";
            when 143 => data_i <= X"033D";
            when 144 => data_i <= X"0347";
            when 145 => data_i <= X"0355";
            when 146 => data_i <= X"0359";
            when 147 => data_i <= X"035B";
            when 148 => data_i <= X"035F";
            when 149 => data_i <= X"036D";
            when 150 => data_i <= X"0371";
            when 151 => data_i <= X"0373";
            when 152 => data_i <= X"0377";
            when 153 => data_i <= X"038B";
            when 154 => data_i <= X"038F";
            when 155 => data_i <= X"0397";
            when 156 => data_i <= X"03A1";
            when 157 => data_i <= X"03A9";
            when 158 => data_i <= X"03AD";
            when 159 => data_i <= X"03B3";
            when 160 => data_i <= X"03B9";
            when 161 => data_i <= X"03C7";
            when 162 => data_i <= X"03CB";
            when 163 => data_i <= X"03D1";
            when 164 => data_i <= X"03D7";
            when 165 => data_i <= X"03DF";
            when 166 => data_i <= X"03E5";
            when 167 => data_i <= X"03F1";
            when 168 => data_i <= X"03F5";
            when 169 => data_i <= X"03FB";
            when 170 => data_i <= X"03FD";
            when 171 => data_i <= X"0407";
            when 172 => data_i <= X"0409";
            when 173 => data_i <= X"040F";
            when 174 => data_i <= X"0419";
            when 175 => data_i <= X"041B";
            when 176 => data_i <= X"0425";
            when 177 => data_i <= X"0427";
            when 178 => data_i <= X"042D";
            when 179 => data_i <= X"043F";
            when 180 => data_i <= X"0443";
            when 181 => data_i <= X"0445";
            when 182 => data_i <= X"0449";
            when 183 => data_i <= X"044F";
            when 184 => data_i <= X"0455";
            when 185 => data_i <= X"045D";
            when 186 => data_i <= X"0463";
            when 187 => data_i <= X"0469";
            when 188 => data_i <= X"047F";
            when 189 => data_i <= X"0481";
            when 190 => data_i <= X"048B";
            when 191 => data_i <= X"0493";
            when 192 => data_i <= X"049D";
            when 193 => data_i <= X"04A3";
            when 194 => data_i <= X"04A9";
            when 195 => data_i <= X"04B1";
            when 196 => data_i <= X"04BD";
            when 197 => data_i <= X"04C1";
            when 198 => data_i <= X"04C7";
            when 199 => data_i <= X"04CD";
            when 200 => data_i <= X"04CF";
            when 201 => data_i <= X"04D5";
            when 202 => data_i <= X"04E1";
            when 203 => data_i <= X"04EB";
            when 204 => data_i <= X"04FD";
            when 205 => data_i <= X"04FF";
            when 206 => data_i <= X"0503";
            when 207 => data_i <= X"0509";
            when 208 => data_i <= X"050B";
            when 209 => data_i <= X"0511";
            when 210 => data_i <= X"0515";
            when 211 => data_i <= X"0517";
            when 212 => data_i <= X"051B";
            when 213 => data_i <= X"0527";
            when 214 => data_i <= X"0529";
            when 215 => data_i <= X"052F";
            when 216 => data_i <= X"0551";
            when 217 => data_i <= X"0557";
            when 218 => data_i <= X"055D";
            when 219 => data_i <= X"0565";
            when 220 => data_i <= X"0577";
            when 221 => data_i <= X"0581";
            when 222 => data_i <= X"058F";
            when 223 => data_i <= X"0593";
            when 224 => data_i <= X"0595";
            when 225 => data_i <= X"0599";
            when 226 => data_i <= X"059F";
            when 227 => data_i <= X"05A7";
            when 228 => data_i <= X"05AB";
            when 229 => data_i <= X"05AD";
            when 230 => data_i <= X"05B3";
            when 231 => data_i <= X"05BF";
            when 232 => data_i <= X"05C9";
            when 233 => data_i <= X"05CB";
            when 234 => data_i <= X"05CF";
            when 235 => data_i <= X"05D1";
            when 236 => data_i <= X"05D5";
            when 237 => data_i <= X"05DB";
            when 238 => data_i <= X"05E7";
            when 239 => data_i <= X"05F3";
            when 240 => data_i <= X"05FB";
            when 241 => data_i <= X"0607";
            when 242 => data_i <= X"060D";
            when 243 => data_i <= X"0611";
            when 244 => data_i <= X"0617";
            when 245 => data_i <= X"061F";
            when 246 => data_i <= X"0623";
            when 247 => data_i <= X"062B";
            when 248 => data_i <= X"062F";
            when 249 => data_i <= X"063D";
            when 250 => data_i <= X"0641";
            when 251 => data_i <= X"0647";
            when 252 => data_i <= X"0649";
            when 253 => data_i <= X"064D";
            when 254 => data_i <= X"0653";
            when 255 => data_i <= X"0655";
            when 256 => data_i <= X"065B";
            when 257 => data_i <= X"0665";
            when 258 => data_i <= X"0679";
            when 259 => data_i <= X"067F";
            when 260 => data_i <= X"0683";
            when 261 => data_i <= X"0685";
            when 262 => data_i <= X"069D";
            when 263 => data_i <= X"06A1";
            when 264 => data_i <= X"06A3";
            when 265 => data_i <= X"06AD";
            when 266 => data_i <= X"06B9";
            when 267 => data_i <= X"06BB";
            when 268 => data_i <= X"06C5";
            when 269 => data_i <= X"06CD";
            when 270 => data_i <= X"06D3";
            when 271 => data_i <= X"06D9";
            when 272 => data_i <= X"06DF";
            when 273 => data_i <= X"06F1";
            when 274 => data_i <= X"06F7";
            when 275 => data_i <= X"06FB";
            when 276 => data_i <= X"06FD";
            when 277 => data_i <= X"0709";
            when 278 => data_i <= X"0713";
            when 279 => data_i <= X"071F";
            when 280 => data_i <= X"0727";
            when 281 => data_i <= X"0737";
            when 282 => data_i <= X"0745";
            when 283 => data_i <= X"074B";
            when 284 => data_i <= X"074F";
            when 285 => data_i <= X"0751";
            when 286 => data_i <= X"0755";
            when 287 => data_i <= X"0757";
            when 288 => data_i <= X"0761";
            when 289 => data_i <= X"076D";
            when 290 => data_i <= X"0773";
            when 291 => data_i <= X"0779";
            when 292 => data_i <= X"078B";
            when 293 => data_i <= X"078D";
            when 294 => data_i <= X"079D";
            when 295 => data_i <= X"079F";
            when 296 => data_i <= X"07B5";
            when 297 => data_i <= X"07BB";
            when 298 => data_i <= X"07C3";
            when 299 => data_i <= X"07C9";
            when 300 => data_i <= X"07CD";
            when 301 => data_i <= X"07CF";
            when 302 => data_i <= X"07D3";
            when 303 => data_i <= X"07DB";
            when 304 => data_i <= X"07E1";
            when 305 => data_i <= X"07EB";
            when 306 => data_i <= X"07ED";
            when 307 => data_i <= X"07F7";
            when 308 => data_i <= X"0805";
            when 309 => data_i <= X"080F";
            when 310 => data_i <= X"0815";
            when 311 => data_i <= X"0821";
            when 312 => data_i <= X"0823";
            when 313 => data_i <= X"0827";
            when 314 => data_i <= X"0829";
            when 315 => data_i <= X"0833";
            when 316 => data_i <= X"083F";
            when 317 => data_i <= X"0841";
            when 318 => data_i <= X"0851";
            when 319 => data_i <= X"0853";
            when 320 => data_i <= X"0859";
            when 321 => data_i <= X"085D";
            when 322 => data_i <= X"085F";
            when 323 => data_i <= X"0869";
            when 324 => data_i <= X"0871";
            when 325 => data_i <= X"0883";
            when 326 => data_i <= X"089B";
            when 327 => data_i <= X"089F";
            when 328 => data_i <= X"08A5";
            when 329 => data_i <= X"08AD";
            when 330 => data_i <= X"08BD";
            when 331 => data_i <= X"08BF";
            when 332 => data_i <= X"08C3";
            when 333 => data_i <= X"08CB";
            when 334 => data_i <= X"08DB";
            when 335 => data_i <= X"08DD";
            when 336 => data_i <= X"08E1";
            when 337 => data_i <= X"08E9";
            when 338 => data_i <= X"08EF";
            when 339 => data_i <= X"08F5";
            when 340 => data_i <= X"08F9";
            when 341 => data_i <= X"0905";
            when 342 => data_i <= X"0907";
            when 343 => data_i <= X"091D";
            when 344 => data_i <= X"0923";
            when 345 => data_i <= X"0925";
            when 346 => data_i <= X"092B";
            when 347 => data_i <= X"092F";
            when 348 => data_i <= X"0935";
            when 349 => data_i <= X"0943";
            when 350 => data_i <= X"0949";
            when 351 => data_i <= X"094D";
            when 352 => data_i <= X"094F";
            when 353 => data_i <= X"0955";
            when 354 => data_i <= X"0959";
            when 355 => data_i <= X"095F";
            when 356 => data_i <= X"096B";
            when 357 => data_i <= X"0971";
            when 358 => data_i <= X"0977";
            when 359 => data_i <= X"0985";
            when 360 => data_i <= X"0989";
            when 361 => data_i <= X"098F";
            when 362 => data_i <= X"099B";
            when 363 => data_i <= X"09A3";
            when 364 => data_i <= X"09A9";
            when 365 => data_i <= X"09AD";
            when 366 => data_i <= X"09C7";
            when 367 => data_i <= X"09D9";
            when 368 => data_i <= X"09E3";
            when 369 => data_i <= X"09EB";
            when 370 => data_i <= X"09EF";
            when 371 => data_i <= X"09F5";
            when 372 => data_i <= X"09F7";
            when 373 => data_i <= X"09FD";
            when 374 => data_i <= X"0A13";
            when 375 => data_i <= X"0A1F";
            when 376 => data_i <= X"0A21";
            when 377 => data_i <= X"0A31";
            when 378 => data_i <= X"0A39";
            when 379 => data_i <= X"0A3D";
            when 380 => data_i <= X"0A49";
            when 381 => data_i <= X"0A57";
            when 382 => data_i <= X"0A61";
            when 383 => data_i <= X"0A63";
            when 384 => data_i <= X"0A67";
            when 385 => data_i <= X"0A6F";
            when 386 => data_i <= X"0A75";
            when 387 => data_i <= X"0A7B";
            when 388 => data_i <= X"0A7F";
            when 389 => data_i <= X"0A81";
            when 390 => data_i <= X"0A85";
            when 391 => data_i <= X"0A8B";
            when 392 => data_i <= X"0A93";
            when 393 => data_i <= X"0A97";
            when 394 => data_i <= X"0A99";
            when 395 => data_i <= X"0A9F";
            when 396 => data_i <= X"0AA9";
            when 397 => data_i <= X"0AAB";
            when 398 => data_i <= X"0AB5";
            when 399 => data_i <= X"0ABD";
            when 400 => data_i <= X"0AC1";
            when 401 => data_i <= X"0ACF";
            when 402 => data_i <= X"0AD9";
            when 403 => data_i <= X"0AE5";
            when 404 => data_i <= X"0AE7";
            when 405 => data_i <= X"0AED";
            when 406 => data_i <= X"0AF1";
            when 407 => data_i <= X"0AF3";
            when 408 => data_i <= X"0B03";
            when 409 => data_i <= X"0B11";
            when 410 => data_i <= X"0B15";
            when 411 => data_i <= X"0B1B";
            when 412 => data_i <= X"0B23";
            when 413 => data_i <= X"0B29";
            when 414 => data_i <= X"0B2D";
            when 415 => data_i <= X"0B3F";
            when 416 => data_i <= X"0B47";
            when 417 => data_i <= X"0B51";
            when 418 => data_i <= X"0B57";
            when 419 => data_i <= X"0B5D";
            when 420 => data_i <= X"0B65";
            when 421 => data_i <= X"0B6F";
            when 422 => data_i <= X"0B7B";
            when 423 => data_i <= X"0B89";
            when 424 => data_i <= X"0B8D";
            when 425 => data_i <= X"0B93";
            when 426 => data_i <= X"0B99";
            when 427 => data_i <= X"0B9B";
            when 428 => data_i <= X"0BB7";
            when 429 => data_i <= X"0BB9";
            when 430 => data_i <= X"0BC3";
            when 431 => data_i <= X"0BCB";
            when 432 => data_i <= X"0BCF";
            when 433 => data_i <= X"0BDD";
            when 434 => data_i <= X"0BE1";
            when 435 => data_i <= X"0BE9";
            when 436 => data_i <= X"0BF5";
            when 437 => data_i <= X"0BFB";
            when 438 => data_i <= X"0C07";
            when 439 => data_i <= X"0C0B";
            when 440 => data_i <= X"0C11";
            when 441 => data_i <= X"0C25";
            when 442 => data_i <= X"0C2F";
            when 443 => data_i <= X"0C31";
            when 444 => data_i <= X"0C41";
            when 445 => data_i <= X"0C5B";
            when 446 => data_i <= X"0C5F";
            when 447 => data_i <= X"0C61";
            when 448 => data_i <= X"0C6D";
            when 449 => data_i <= X"0C73";
            when 450 => data_i <= X"0C77";
            when 451 => data_i <= X"0C83";
            when 452 => data_i <= X"0C89";
            when 453 => data_i <= X"0C91";
            when 454 => data_i <= X"0C95";
            when 455 => data_i <= X"0C9D";
            when 456 => data_i <= X"0CB3";
            when 457 => data_i <= X"0CB5";
            when 458 => data_i <= X"0CB9";
            when 459 => data_i <= X"0CBB";
            when 460 => data_i <= X"0CC7";
            when 461 => data_i <= X"0CE3";
            when 462 => data_i <= X"0CE5";
            when 463 => data_i <= X"0CEB";
            when 464 => data_i <= X"0CF1";
            when 465 => data_i <= X"0CF7";
            when 466 => data_i <= X"0CFB";
            when 467 => data_i <= X"0D01";
            when 468 => data_i <= X"0D03";
            when 469 => data_i <= X"0D0F";
            when 470 => data_i <= X"0D13";
            when 471 => data_i <= X"0D1F";
            when 472 => data_i <= X"0D21";
            when 473 => data_i <= X"0D2B";
            when 474 => data_i <= X"0D2D";
            when 475 => data_i <= X"0D3D";
            when 476 => data_i <= X"0D3F";
            when 477 => data_i <= X"0D4F";
            when 478 => data_i <= X"0D55";
            when 479 => data_i <= X"0D69";
            when 480 => data_i <= X"0D79";
            when 481 => data_i <= X"0D81";
            when 482 => data_i <= X"0D85";
            when 483 => data_i <= X"0D87";
            when 484 => data_i <= X"0D8B";
            when 485 => data_i <= X"0D8D";
            when 486 => data_i <= X"0DA3";
            when 487 => data_i <= X"0DAB";
            when 488 => data_i <= X"0DB7";
            when 489 => data_i <= X"0DBD";
            when 490 => data_i <= X"0DC7";
            when 491 => data_i <= X"0DC9";
            when 492 => data_i <= X"0DCD";
            when 493 => data_i <= X"0DD3";
            when 494 => data_i <= X"0DD5";
            when 495 => data_i <= X"0DDB";
            when 496 => data_i <= X"0DE5";
            when 497 => data_i <= X"0DE7";
            when 498 => data_i <= X"0DF3";
            when 499 => data_i <= X"0DFD";
            when 500 => data_i <= X"0DFF";
            when 501 => data_i <= X"0E09";
            when 502 => data_i <= X"0E17";
            when 503 => data_i <= X"0E1D";
            when 504 => data_i <= X"0E21";
            when 505 => data_i <= X"0E27";
            when 506 => data_i <= X"0E2F";
            when 507 => data_i <= X"0E35";
            when 508 => data_i <= X"0E3B";
            when 509 => data_i <= X"0E4B";
            when 510 => data_i <= X"0E57";
            when 511 => data_i <= X"0E59";
            when 512 => data_i <= X"0E5D";
            when 513 => data_i <= X"0E6B";
            when 514 => data_i <= X"0E71";
            when 515 => data_i <= X"0E75";
            when 516 => data_i <= X"0E7D";
            when 517 => data_i <= X"0E87";
            when 518 => data_i <= X"0E8F";
            when 519 => data_i <= X"0E95";
            when 520 => data_i <= X"0E9B";
            when 521 => data_i <= X"0EB1";
            when 522 => data_i <= X"0EB7";
            when 523 => data_i <= X"0EB9";
            when 524 => data_i <= X"0EC3";
            when 525 => data_i <= X"0ED1";
            when 526 => data_i <= X"0ED5";
            when 527 => data_i <= X"0EDB";
            when 528 => data_i <= X"0EED";
            when 529 => data_i <= X"0EEF";
            when 530 => data_i <= X"0EF9";
            when 531 => data_i <= X"0F07";
            when 532 => data_i <= X"0F0B";
            when 533 => data_i <= X"0F0D";
            when 534 => data_i <= X"0F17";
            when 535 => data_i <= X"0F25";
            when 536 => data_i <= X"0F29";
            when 537 => data_i <= X"0F31";
            when 538 => data_i <= X"0F43";
            when 539 => data_i <= X"0F47";
            when 540 => data_i <= X"0F4D";
            when 541 => data_i <= X"0F4F";
            when 542 => data_i <= X"0F53";
            when 543 => data_i <= X"0F59";
            when 544 => data_i <= X"0F5B";
            when 545 => data_i <= X"0F67";
            when 546 => data_i <= X"0F6B";
            when 547 => data_i <= X"0F7F";
            when 548 => data_i <= X"0F95";
            when 549 => data_i <= X"0FA1";
            when 550 => data_i <= X"0FA3";
            when 551 => data_i <= X"0FA7";
            when 552 => data_i <= X"0FAD";
            when 553 => data_i <= X"0FB3";
            when 554 => data_i <= X"0FB5";
            when 555 => data_i <= X"0FBB";
            when 556 => data_i <= X"0FD1";
            when 557 => data_i <= X"0FD3";
            when 558 => data_i <= X"0FD9";
            when 559 => data_i <= X"0FE9";
            when 560 => data_i <= X"0FEF";
            when 561 => data_i <= X"0FFB";
            when 562 => data_i <= X"0FFD";
            when 563 => data_i <= X"1003";
            when 564 => data_i <= X"100F";
            when 565 => data_i <= X"101F";
            when 566 => data_i <= X"1021";
            when 567 => data_i <= X"1025";
            when 568 => data_i <= X"102B";
            when 569 => data_i <= X"1039";
            when 570 => data_i <= X"103D";
            when 571 => data_i <= X"103F";
            when 572 => data_i <= X"1051";
            when 573 => data_i <= X"1069";
            when 574 => data_i <= X"1073";
            when 575 => data_i <= X"1079";
            when 576 => data_i <= X"107B";
            when 577 => data_i <= X"1085";
            when 578 => data_i <= X"1087";
            when 579 => data_i <= X"1091";
            when 580 => data_i <= X"1093";
            when 581 => data_i <= X"109D";
            when 582 => data_i <= X"10A3";
            when 583 => data_i <= X"10A5";
            when 584 => data_i <= X"10AF";
            when 585 => data_i <= X"10B1";
            when 586 => data_i <= X"10BB";
            when 587 => data_i <= X"10C1";
            when 588 => data_i <= X"10C9";
            when 589 => data_i <= X"10E7";
            when 590 => data_i <= X"10F1";
            when 591 => data_i <= X"10F3";
            when 592 => data_i <= X"10FD";
            when 593 => data_i <= X"1105";
            when 594 => data_i <= X"110B";
            when 595 => data_i <= X"1115";
            when 596 => data_i <= X"1127";
            when 597 => data_i <= X"112D";
            when 598 => data_i <= X"1139";
            when 599 => data_i <= X"1145";
            when 600 => data_i <= X"1147";
            when 601 => data_i <= X"1159";
            when 602 => data_i <= X"115F";
            when 603 => data_i <= X"1163";
            when 604 => data_i <= X"1169";
            when 605 => data_i <= X"116F";
            when 606 => data_i <= X"1181";
            when 607 => data_i <= X"1183";
            when 608 => data_i <= X"118D";
            when 609 => data_i <= X"119B";
            when 610 => data_i <= X"11A1";
            when 611 => data_i <= X"11A5";
            when 612 => data_i <= X"11A7";
            when 613 => data_i <= X"11AB";
            when 614 => data_i <= X"11C3";
            when 615 => data_i <= X"11C5";
            when 616 => data_i <= X"11D1";
            when 617 => data_i <= X"11D7";
            when 618 => data_i <= X"11E7";
            when 619 => data_i <= X"11EF";
            when 620 => data_i <= X"11F5";
            when 621 => data_i <= X"11FB";
            when 622 => data_i <= X"120D";
            when 623 => data_i <= X"121D";
            when 624 => data_i <= X"121F";
            when 625 => data_i <= X"1223";
            when 626 => data_i <= X"1229";
            when 627 => data_i <= X"122B";
            when 628 => data_i <= X"1231";
            when 629 => data_i <= X"1237";
            when 630 => data_i <= X"1241";
            when 631 => data_i <= X"1247";
            when 632 => data_i <= X"1253";
            when 633 => data_i <= X"125F";
            when 634 => data_i <= X"1271";
            when 635 => data_i <= X"1273";
            when 636 => data_i <= X"1279";
            when 637 => data_i <= X"127D";
            when 638 => data_i <= X"128F";
            when 639 => data_i <= X"1297";
            when 640 => data_i <= X"12AF";
            when 641 => data_i <= X"12B3";
            when 642 => data_i <= X"12B5";
            when 643 => data_i <= X"12B9";
            when 644 => data_i <= X"12BF";
            when 645 => data_i <= X"12C1";
            when 646 => data_i <= X"12CD";
            when 647 => data_i <= X"12D1";
            when 648 => data_i <= X"12DF";
            when 649 => data_i <= X"12FD";
            when 650 => data_i <= X"1307";
            when 651 => data_i <= X"130D";
            when 652 => data_i <= X"1319";
            when 653 => data_i <= X"1327";
            when 654 => data_i <= X"132D";
            when 655 => data_i <= X"1337";
            when 656 => data_i <= X"1343";
            when 657 => data_i <= X"1345";
            when 658 => data_i <= X"1349";
            when 659 => data_i <= X"134F";
            when 660 => data_i <= X"1357";
            when 661 => data_i <= X"135D";
            when 662 => data_i <= X"1367";
            when 663 => data_i <= X"1369";
            when 664 => data_i <= X"136D";
            when 665 => data_i <= X"137B";
            when 666 => data_i <= X"1381";
            when 667 => data_i <= X"1387";
            when 668 => data_i <= X"138B";
            when 669 => data_i <= X"1391";
            when 670 => data_i <= X"1393";
            when 671 => data_i <= X"139D";
            when 672 => data_i <= X"139F";
            when 673 => data_i <= X"13AF";
            when 674 => data_i <= X"13BB";
            when 675 => data_i <= X"13C3";
            when 676 => data_i <= X"13D5";
            when 677 => data_i <= X"13D9";
            when 678 => data_i <= X"13DF";
            when 679 => data_i <= X"13EB";
            when 680 => data_i <= X"13ED";
            when 681 => data_i <= X"13F3";
            when 682 => data_i <= X"13F9";
            when 683 => data_i <= X"13FF";
            when 684 => data_i <= X"141B";
            when 685 => data_i <= X"1421";
            when 686 => data_i <= X"142F";
            when 687 => data_i <= X"1433";
            when 688 => data_i <= X"143B";
            when 689 => data_i <= X"1445";
            when 690 => data_i <= X"144D";
            when 691 => data_i <= X"1459";
            when 692 => data_i <= X"146B";
            when 693 => data_i <= X"146F";
            when 694 => data_i <= X"1471";
            when 695 => data_i <= X"1475";
            when 696 => data_i <= X"148D";
            when 697 => data_i <= X"1499";
            when 698 => data_i <= X"149F";
            when 699 => data_i <= X"14A1";
            when 700 => data_i <= X"14B1";
            when 701 => data_i <= X"14B7";
            when 702 => data_i <= X"14BD";
            when 703 => data_i <= X"14CB";
            when 704 => data_i <= X"14D5";
            when 705 => data_i <= X"14E3";
            when 706 => data_i <= X"14E7";
            when 707 => data_i <= X"1505";
            when 708 => data_i <= X"150B";
            when 709 => data_i <= X"1511";
            when 710 => data_i <= X"1517";
            when 711 => data_i <= X"151F";
            when 712 => data_i <= X"1525";
            when 713 => data_i <= X"1529";
            when 714 => data_i <= X"152B";
            when 715 => data_i <= X"1537";
            when 716 => data_i <= X"153D";
            when 717 => data_i <= X"1541";
            when 718 => data_i <= X"1543";
            when 719 => data_i <= X"1549";
            when 720 => data_i <= X"155F";
            when 721 => data_i <= X"1565";
            when 722 => data_i <= X"1567";
            when 723 => data_i <= X"156B";
            when 724 => data_i <= X"157D";
            when 725 => data_i <= X"157F";
            when 726 => data_i <= X"1583";
            when 727 => data_i <= X"158F";
            when 728 => data_i <= X"1591";
            when 729 => data_i <= X"1597";
            when 730 => data_i <= X"159B";
            when 731 => data_i <= X"15B5";
            when 732 => data_i <= X"15BB";
            when 733 => data_i <= X"15C1";
            when 734 => data_i <= X"15C5";
            when 735 => data_i <= X"15CD";
            when 736 => data_i <= X"15D7";
            when 737 => data_i <= X"15F7";
            when 738 => data_i <= X"1607";
            when 739 => data_i <= X"1609";
            when 740 => data_i <= X"160F";
            when 741 => data_i <= X"1613";
            when 742 => data_i <= X"1615";
            when 743 => data_i <= X"1619";
            when 744 => data_i <= X"161B";
            when 745 => data_i <= X"1625";
            when 746 => data_i <= X"1633";
            when 747 => data_i <= X"1639";
            when 748 => data_i <= X"163D";
            when 749 => data_i <= X"1645";
            when 750 => data_i <= X"164F";
            when 751 => data_i <= X"1655";
            when 752 => data_i <= X"1669";
            when 753 => data_i <= X"166D";
            when 754 => data_i <= X"166F";
            when 755 => data_i <= X"1675";
            when 756 => data_i <= X"1693";
            when 757 => data_i <= X"1697";
            when 758 => data_i <= X"169F";
            when 759 => data_i <= X"16A9";
            when 760 => data_i <= X"16AF";
            when 761 => data_i <= X"16B5";
            when 762 => data_i <= X"16BD";
            when 763 => data_i <= X"16C3";
            when 764 => data_i <= X"16CF";
            when 765 => data_i <= X"16D3";
            when 766 => data_i <= X"16D9";
            when 767 => data_i <= X"16DB";
            when 768 => data_i <= X"16E1";
            when 769 => data_i <= X"16E5";
            when 770 => data_i <= X"16EB";
            when 771 => data_i <= X"16ED";
            when 772 => data_i <= X"16F7";
            when 773 => data_i <= X"16F9";
            when 774 => data_i <= X"1709";
            when 775 => data_i <= X"170F";
            when 776 => data_i <= X"1723";
            when 777 => data_i <= X"1727";
            when 778 => data_i <= X"1733";
            when 779 => data_i <= X"1741";
            when 780 => data_i <= X"175D";
            when 781 => data_i <= X"1763";
            when 782 => data_i <= X"1777";
            when 783 => data_i <= X"177B";
            when 784 => data_i <= X"178D";
            when 785 => data_i <= X"1795";
            when 786 => data_i <= X"179B";
            when 787 => data_i <= X"179F";
            when 788 => data_i <= X"17A5";
            when 789 => data_i <= X"17B3";
            when 790 => data_i <= X"17B9";
            when 791 => data_i <= X"17BF";
            when 792 => data_i <= X"17C9";
            when 793 => data_i <= X"17CB";
            when 794 => data_i <= X"17D5";
            when 795 => data_i <= X"17E1";
            when 796 => data_i <= X"17E9";
            when 797 => data_i <= X"17F3";
            when 798 => data_i <= X"17F5";
            when 799 => data_i <= X"17FF";
            when 800 => data_i <= X"1807";
            when 801 => data_i <= X"1813";
            when 802 => data_i <= X"181D";
            when 803 => data_i <= X"1835";
            when 804 => data_i <= X"1837";
            when 805 => data_i <= X"183B";
            when 806 => data_i <= X"1843";
            when 807 => data_i <= X"1849";
            when 808 => data_i <= X"184D";
            when 809 => data_i <= X"1855";
            when 810 => data_i <= X"1867";
            when 811 => data_i <= X"1871";
            when 812 => data_i <= X"1877";
            when 813 => data_i <= X"187D";
            when 814 => data_i <= X"187F";
            when 815 => data_i <= X"1885";
            when 816 => data_i <= X"188F";
            when 817 => data_i <= X"189B";
            when 818 => data_i <= X"189D";
            when 819 => data_i <= X"18A7";
            when 820 => data_i <= X"18AD";
            when 821 => data_i <= X"18B3";
            when 822 => data_i <= X"18B9";
            when 823 => data_i <= X"18C1";
            when 824 => data_i <= X"18C7";
            when 825 => data_i <= X"18D1";
            when 826 => data_i <= X"18D7";
            when 827 => data_i <= X"18D9";
            when 828 => data_i <= X"18DF";
            when 829 => data_i <= X"18E5";
            when 830 => data_i <= X"18EB";
            when 831 => data_i <= X"18F5";
            when 832 => data_i <= X"18FD";
            when 833 => data_i <= X"1915";
            when 834 => data_i <= X"191B";
            when 835 => data_i <= X"1931";
            when 836 => data_i <= X"1933";
            when 837 => data_i <= X"1945";
            when 838 => data_i <= X"1949";
            when 839 => data_i <= X"1951";
            when 840 => data_i <= X"195B";
            when 841 => data_i <= X"1979";
            when 842 => data_i <= X"1981";
            when 843 => data_i <= X"1993";
            when 844 => data_i <= X"1997";
            when 845 => data_i <= X"1999";
            when 846 => data_i <= X"19A3";
            when 847 => data_i <= X"19A9";
            when 848 => data_i <= X"19AB";
            when 849 => data_i <= X"19B1";
            when 850 => data_i <= X"19B5";
            when 851 => data_i <= X"19C7";
            when 852 => data_i <= X"19CF";
            when 853 => data_i <= X"19DB";
            when 854 => data_i <= X"19ED";
            when 855 => data_i <= X"19FD";
            when 856 => data_i <= X"1A03";
            when 857 => data_i <= X"1A05";
            when 858 => data_i <= X"1A11";
            when 859 => data_i <= X"1A17";
            when 860 => data_i <= X"1A21";
            when 861 => data_i <= X"1A23";
            when 862 => data_i <= X"1A2D";
            when 863 => data_i <= X"1A2F";
            when 864 => data_i <= X"1A35";
            when 865 => data_i <= X"1A3F";
            when 866 => data_i <= X"1A4D";
            when 867 => data_i <= X"1A51";
            when 868 => data_i <= X"1A69";
            when 869 => data_i <= X"1A6B";
            when 870 => data_i <= X"1A7B";
            when 871 => data_i <= X"1A7D";
            when 872 => data_i <= X"1A87";
            when 873 => data_i <= X"1A89";
            when 874 => data_i <= X"1A93";
            when 875 => data_i <= X"1AA7";
            when 876 => data_i <= X"1AAB";
            when 877 => data_i <= X"1AAD";
            when 878 => data_i <= X"1AB1";
            when 879 => data_i <= X"1AB9";
            when 880 => data_i <= X"1AC9";
            when 881 => data_i <= X"1ACF";
            when 882 => data_i <= X"1AD5";
            when 883 => data_i <= X"1AD7";
            when 884 => data_i <= X"1AE3";
            when 885 => data_i <= X"1AF3";
            when 886 => data_i <= X"1AFB";
            when 887 => data_i <= X"1AFF";
            when 888 => data_i <= X"1B05";
            when 889 => data_i <= X"1B23";
            when 890 => data_i <= X"1B25";
            when 891 => data_i <= X"1B2F";
            when 892 => data_i <= X"1B31";
            when 893 => data_i <= X"1B37";
            when 894 => data_i <= X"1B3B";
            when 895 => data_i <= X"1B41";
            when 896 => data_i <= X"1B47";
            when 897 => data_i <= X"1B4F";
            when 898 => data_i <= X"1B55";
            when 899 => data_i <= X"1B59";
            when 900 => data_i <= X"1B65";
            when 901 => data_i <= X"1B6B";
            when 902 => data_i <= X"1B73";
            when 903 => data_i <= X"1B7F";
            when 904 => data_i <= X"1B83";
            when 905 => data_i <= X"1B91";
            when 906 => data_i <= X"1B9D";
            when 907 => data_i <= X"1BA7";
            when 908 => data_i <= X"1BBF";
            when 909 => data_i <= X"1BC5";
            when 910 => data_i <= X"1BD1";
            when 911 => data_i <= X"1BD7";
            when 912 => data_i <= X"1BD9";
            when 913 => data_i <= X"1BEF";
            when 914 => data_i <= X"1BF7";
            when 915 => data_i <= X"1C09";
            when 916 => data_i <= X"1C13";
            when 917 => data_i <= X"1C19";
            when 918 => data_i <= X"1C27";
            when 919 => data_i <= X"1C2B";
            when 920 => data_i <= X"1C2D";
            when 921 => data_i <= X"1C33";
            when 922 => data_i <= X"1C3D";
            when 923 => data_i <= X"1C45";
            when 924 => data_i <= X"1C4B";
            when 925 => data_i <= X"1C4F";
            when 926 => data_i <= X"1C55";
            when 927 => data_i <= X"1C73";
            when 928 => data_i <= X"1C81";
            when 929 => data_i <= X"1C8B";
            when 930 => data_i <= X"1C8D";
            when 931 => data_i <= X"1C99";
            when 932 => data_i <= X"1CA3";
            when 933 => data_i <= X"1CA5";
            when 934 => data_i <= X"1CB5";
            when 935 => data_i <= X"1CB7";
            when 936 => data_i <= X"1CC9";
            when 937 => data_i <= X"1CE1";
            when 938 => data_i <= X"1CF3";
            when 939 => data_i <= X"1CF9";
            when 940 => data_i <= X"1D09";
            when 941 => data_i <= X"1D1B";
            when 942 => data_i <= X"1D21";
            when 943 => data_i <= X"1D23";
            when 944 => data_i <= X"1D35";
            when 945 => data_i <= X"1D39";
            when 946 => data_i <= X"1D3F";
            when 947 => data_i <= X"1D41";
            when 948 => data_i <= X"1D4B";
            when 949 => data_i <= X"1D53";
            when 950 => data_i <= X"1D5D";
            when 951 => data_i <= X"1D63";
            when 952 => data_i <= X"1D69";
            when 953 => data_i <= X"1D71";
            when 954 => data_i <= X"1D75";
            when 955 => data_i <= X"1D7B";
            when 956 => data_i <= X"1D7D";
            when 957 => data_i <= X"1D87";
            when 958 => data_i <= X"1D89";
            when 959 => data_i <= X"1D95";
            when 960 => data_i <= X"1D99";
            when 961 => data_i <= X"1D9F";
            when 962 => data_i <= X"1DA5";
            when 963 => data_i <= X"1DA7";
            when 964 => data_i <= X"1DB3";
            when 965 => data_i <= X"1DB7";
            when 966 => data_i <= X"1DC5";
            when 967 => data_i <= X"1DD7";
            when 968 => data_i <= X"1DDB";
            when 969 => data_i <= X"1DE1";
            when 970 => data_i <= X"1DF5";
            when 971 => data_i <= X"1DF9";
            when 972 => data_i <= X"1E01";
            when 973 => data_i <= X"1E07";
            when 974 => data_i <= X"1E0B";
            when 975 => data_i <= X"1E13";
            when 976 => data_i <= X"1E17";
            when 977 => data_i <= X"1E25";
            when 978 => data_i <= X"1E2B";
            when 979 => data_i <= X"1E2F";
            when 980 => data_i <= X"1E3D";
            when 981 => data_i <= X"1E49";
            when 982 => data_i <= X"1E4D";
            when 983 => data_i <= X"1E4F";
            when 984 => data_i <= X"1E6D";
            when 985 => data_i <= X"1E71";
            when 986 => data_i <= X"1E89";
            when 987 => data_i <= X"1E8F";
            when 988 => data_i <= X"1E95";
            when 989 => data_i <= X"1EA1";
            when 990 => data_i <= X"1EAD";
            when 991 => data_i <= X"1EBB";
            when 992 => data_i <= X"1EC1";
            when 993 => data_i <= X"1EC5";
            when 994 => data_i <= X"1EC7";
            when 995 => data_i <= X"1ECB";
            when 996 => data_i <= X"1EDD";
            when 997 => data_i <= X"1EE3";
            when 998 => data_i <= X"1EEF";
            when 999 => data_i <= X"1EF7";
            when 1000 => data_i <= X"1EFD";
            when 1001 => data_i <= X"1F01";
            when 1002 => data_i <= X"1F0D";
            when 1003 => data_i <= X"1F0F";
            when 1004 => data_i <= X"1F1B";
            when 1005 => data_i <= X"1F39";
            when 1006 => data_i <= X"1F49";
            when 1007 => data_i <= X"1F4B";
            when 1008 => data_i <= X"1F51";
            when 1009 => data_i <= X"1F67";
            when 1010 => data_i <= X"1F75";
            when 1011 => data_i <= X"1F7B";
            when 1012 => data_i <= X"1F85";
            when 1013 => data_i <= X"1F91";
            when 1014 => data_i <= X"1F97";
            when 1015 => data_i <= X"1F99";
            when 1016 => data_i <= X"1F9D";
            when 1017 => data_i <= X"1FA5";
            when 1018 => data_i <= X"1FAF";
            when 1019 => data_i <= X"1FB5";
            when 1020 => data_i <= X"1FBB";
            when 1021 => data_i <= X"1FD3";
            when 1022 => data_i <= X"1FE1";
            when 1023 => data_i <= X"1FE7";
            when 1024 => data_i <= X"1FEB";
            when 1025 => data_i <= X"1FF3";
            when 1026 => data_i <= X"1FFF";
            when 1027 => data_i <= X"2011";
            when 1028 => data_i <= X"201B";
            when 1029 => data_i <= X"201D";
            when 1030 => data_i <= X"2027";
            when 1031 => data_i <= X"2029";
            when 1032 => data_i <= X"202D";
            when 1033 => data_i <= X"2033";
            when 1034 => data_i <= X"2047";
            when 1035 => data_i <= X"204D";
            when 1036 => data_i <= X"2051";
            when 1037 => data_i <= X"205F";
            when 1038 => data_i <= X"2063";
            when 1039 => data_i <= X"2065";
            when 1040 => data_i <= X"2069";
            when 1041 => data_i <= X"2077";
            when 1042 => data_i <= X"207D";
            when 1043 => data_i <= X"2089";
            when 1044 => data_i <= X"20A1";
            when 1045 => data_i <= X"20AB";
            when 1046 => data_i <= X"20B1";
            when 1047 => data_i <= X"20B9";
            when 1048 => data_i <= X"20C3";
            when 1049 => data_i <= X"20C5";
            when 1050 => data_i <= X"20E3";
            when 1051 => data_i <= X"20E7";
            when 1052 => data_i <= X"20ED";
            when 1053 => data_i <= X"20EF";
            when 1054 => data_i <= X"20FB";
            when 1055 => data_i <= X"20FF";
            when 1056 => data_i <= X"210D";
            when 1057 => data_i <= X"2113";
            when 1058 => data_i <= X"2135";
            when 1059 => data_i <= X"2141";
            when 1060 => data_i <= X"2149";
            when 1061 => data_i <= X"214F";
            when 1062 => data_i <= X"2159";
            when 1063 => data_i <= X"215B";
            when 1064 => data_i <= X"215F";
            when 1065 => data_i <= X"2173";
            when 1066 => data_i <= X"217D";
            when 1067 => data_i <= X"2185";
            when 1068 => data_i <= X"2195";
            when 1069 => data_i <= X"2197";
            when 1070 => data_i <= X"21A1";
            when 1071 => data_i <= X"21AF";
            when 1072 => data_i <= X"21B3";
            when 1073 => data_i <= X"21B5";
            when 1074 => data_i <= X"21C1";
            when 1075 => data_i <= X"21C7";
            when 1076 => data_i <= X"21D7";
            when 1077 => data_i <= X"21DD";
            when 1078 => data_i <= X"21E5";
            when 1079 => data_i <= X"21E9";
            when 1080 => data_i <= X"21F1";
            when 1081 => data_i <= X"21F5";
            when 1082 => data_i <= X"21FB";
            when 1083 => data_i <= X"2203";
            when 1084 => data_i <= X"2209";
            when 1085 => data_i <= X"220F";
            when 1086 => data_i <= X"221B";
            when 1087 => data_i <= X"2221";
            when 1088 => data_i <= X"2225";
            when 1089 => data_i <= X"222B";
            when 1090 => data_i <= X"2231";
            when 1091 => data_i <= X"2239";
            when 1092 => data_i <= X"224B";
            when 1093 => data_i <= X"224F";
            when 1094 => data_i <= X"2263";
            when 1095 => data_i <= X"2267";
            when 1096 => data_i <= X"2273";
            when 1097 => data_i <= X"2275";
            when 1098 => data_i <= X"227F";
            when 1099 => data_i <= X"2285";
            when 1100 => data_i <= X"2287";
            when 1101 => data_i <= X"2291";
            when 1102 => data_i <= X"229D";
            when 1103 => data_i <= X"229F";
            when 1104 => data_i <= X"22A3";
            when 1105 => data_i <= X"22B7";
            when 1106 => data_i <= X"22BD";
            when 1107 => data_i <= X"22DB";
            when 1108 => data_i <= X"22E1";
            when 1109 => data_i <= X"22E5";
            when 1110 => data_i <= X"22ED";
            when 1111 => data_i <= X"22F7";
            when 1112 => data_i <= X"2303";
            when 1113 => data_i <= X"2309";
            when 1114 => data_i <= X"230B";
            when 1115 => data_i <= X"2327";
            when 1116 => data_i <= X"2329";
            when 1117 => data_i <= X"232F";
            when 1118 => data_i <= X"2333";
            when 1119 => data_i <= X"2335";
            when 1120 => data_i <= X"2345";
            when 1121 => data_i <= X"2351";
            when 1122 => data_i <= X"2353";
            when 1123 => data_i <= X"2359";
            when 1124 => data_i <= X"2363";
            when 1125 => data_i <= X"236B";
            when 1126 => data_i <= X"2383";
            when 1127 => data_i <= X"238F";
            when 1128 => data_i <= X"2395";
            when 1129 => data_i <= X"23A7";
            when 1130 => data_i <= X"23AD";
            when 1131 => data_i <= X"23B1";
            when 1132 => data_i <= X"23BF";
            when 1133 => data_i <= X"23C5";
            when 1134 => data_i <= X"23C9";
            when 1135 => data_i <= X"23D5";
            when 1136 => data_i <= X"23DD";
            when 1137 => data_i <= X"23E3";
            when 1138 => data_i <= X"23EF";
            when 1139 => data_i <= X"23F3";
            when 1140 => data_i <= X"23F9";
            when 1141 => data_i <= X"2405";
            when 1142 => data_i <= X"240B";
            when 1143 => data_i <= X"2417";
            when 1144 => data_i <= X"2419";
            when 1145 => data_i <= X"2429";
            when 1146 => data_i <= X"243D";
            when 1147 => data_i <= X"2441";
            when 1148 => data_i <= X"2443";
            when 1149 => data_i <= X"244D";
            when 1150 => data_i <= X"245F";
            when 1151 => data_i <= X"2467";
            when 1152 => data_i <= X"246B";
            when 1153 => data_i <= X"2479";
            when 1154 => data_i <= X"247D";
            when 1155 => data_i <= X"247F";
            when 1156 => data_i <= X"2485";
            when 1157 => data_i <= X"249B";
            when 1158 => data_i <= X"24A1";
            when 1159 => data_i <= X"24AF";
            when 1160 => data_i <= X"24B5";
            when 1161 => data_i <= X"24BB";
            when 1162 => data_i <= X"24C5";
            when 1163 => data_i <= X"24CB";
            when 1164 => data_i <= X"24CD";
            when 1165 => data_i <= X"24D7";
            when 1166 => data_i <= X"24D9";
            when 1167 => data_i <= X"24DD";
            when 1168 => data_i <= X"24DF";
            when 1169 => data_i <= X"24F5";
            when 1170 => data_i <= X"24F7";
            when 1171 => data_i <= X"24FB";
            when 1172 => data_i <= X"2501";
            when 1173 => data_i <= X"2507";
            when 1174 => data_i <= X"2513";
            when 1175 => data_i <= X"2519";
            when 1176 => data_i <= X"2527";
            when 1177 => data_i <= X"2531";
            when 1178 => data_i <= X"253D";
            when 1179 => data_i <= X"2543";
            when 1180 => data_i <= X"254B";
            when 1181 => data_i <= X"254F";
            when 1182 => data_i <= X"2573";
            when 1183 => data_i <= X"2581";
            when 1184 => data_i <= X"258D";
            when 1185 => data_i <= X"2593";
            when 1186 => data_i <= X"2597";
            when 1187 => data_i <= X"259D";
            when 1188 => data_i <= X"259F";
            when 1189 => data_i <= X"25AB";
            when 1190 => data_i <= X"25B1";
            when 1191 => data_i <= X"25BD";
            when 1192 => data_i <= X"25CD";
            when 1193 => data_i <= X"25CF";
            when 1194 => data_i <= X"25D9";
            when 1195 => data_i <= X"25E1";
            when 1196 => data_i <= X"25F7";
            when 1197 => data_i <= X"25F9";
            when 1198 => data_i <= X"2605";
            when 1199 => data_i <= X"260B";
            when 1200 => data_i <= X"260F";
            when 1201 => data_i <= X"2615";
            when 1202 => data_i <= X"2627";
            when 1203 => data_i <= X"2629";
            when 1204 => data_i <= X"2635";
            when 1205 => data_i <= X"263B";
            when 1206 => data_i <= X"263F";
            when 1207 => data_i <= X"264B";
            when 1208 => data_i <= X"2653";
            when 1209 => data_i <= X"2659";
            when 1210 => data_i <= X"2665";
            when 1211 => data_i <= X"2669";
            when 1212 => data_i <= X"266F";
            when 1213 => data_i <= X"267B";
            when 1214 => data_i <= X"2681";
            when 1215 => data_i <= X"2683";
            when 1216 => data_i <= X"268F";
            when 1217 => data_i <= X"269B";
            when 1218 => data_i <= X"269F";
            when 1219 => data_i <= X"26AD";
            when 1220 => data_i <= X"26B3";
            when 1221 => data_i <= X"26C3";
            when 1222 => data_i <= X"26C9";
            when 1223 => data_i <= X"26CB";
            when 1224 => data_i <= X"26D5";
            when 1225 => data_i <= X"26DD";
            when 1226 => data_i <= X"26EF";
            when 1227 => data_i <= X"26F5";
            when others => data_i <= data_i;
        end case;
    end if;
end process;

DATA <= data_i;


end RTL;    --PRIME_ROM