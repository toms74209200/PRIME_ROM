/* ============================================================================
 *  Title       : Prime number ROM
 *
 *  File Name	: PRIME_ROM.v
 *  Project     :
 *  Block       :
 *  Tree        :
 *  Designer    : toms74209200 <https://github.com/toms74209200>
 *  Created     : 2019/09/22
 *  Copyright   : 2019 toms74209200
 *  License     : MIT License.
 *                http://opensource.org/licenses/mit-license.php
 * ============================================================================*/
module PRIME_ROM
    (
    // System
    CLK,        //(p) Clock

    // ROM interface
    ADDRESS,    //(p) Address
    DATA        //(p) Data
    );

// Port
// System
input           CLK;        //(p) Clock

// ROM interface
input  [10:0]   ADDRESS;    //(p) Address
output [15:0]   DATA;       //(p) Data

// Internal signals
reg [15:0]      rom_prime[0:1227];  // ROM table
reg [15:0]      data_i;             // Data

/* ============================================================================
 * ROM table
 * ============================================================================*/
initial begin
rom_prime[0]    = 16'h0003;
rom_prime[1]    = 16'h0005;
rom_prime[2]    = 16'h0007;
rom_prime[3]    = 16'h000B;
rom_prime[4]    = 16'h000D;
rom_prime[5]    = 16'h0011;
rom_prime[6]    = 16'h0013;
rom_prime[7]    = 16'h0017;
rom_prime[8]    = 16'h001D;
rom_prime[9]    = 16'h001F;
rom_prime[10]   = 16'h0025;
rom_prime[11]   = 16'h0029;
rom_prime[12]   = 16'h002B;
rom_prime[13]   = 16'h002F;
rom_prime[14]   = 16'h0035;
rom_prime[15]   = 16'h003B;
rom_prime[16]   = 16'h003D;
rom_prime[17]   = 16'h0043;
rom_prime[18]   = 16'h0047;
rom_prime[19]   = 16'h0049;
rom_prime[20]   = 16'h004F;
rom_prime[21]   = 16'h0053;
rom_prime[22]   = 16'h0059;
rom_prime[23]   = 16'h0061;
rom_prime[24]   = 16'h0065;
rom_prime[25]   = 16'h0067;
rom_prime[26]   = 16'h006B;
rom_prime[27]   = 16'h006D;
rom_prime[28]   = 16'h0071;
rom_prime[29]   = 16'h007F;
rom_prime[30]   = 16'h0083;
rom_prime[31]   = 16'h0089;
rom_prime[32]   = 16'h008B;
rom_prime[33]   = 16'h0095;
rom_prime[34]   = 16'h0097;
rom_prime[35]   = 16'h009D;
rom_prime[36]   = 16'h00A3;
rom_prime[37]   = 16'h00A7;
rom_prime[38]   = 16'h00AD;
rom_prime[39]   = 16'h00B3;
rom_prime[40]   = 16'h00B5;
rom_prime[41]   = 16'h00BF;
rom_prime[42]   = 16'h00C1;
rom_prime[43]   = 16'h00C5;
rom_prime[44]   = 16'h00C7;
rom_prime[45]   = 16'h00D3;
rom_prime[46]   = 16'h00DF;
rom_prime[47]   = 16'h00E3;
rom_prime[48]   = 16'h00E5;
rom_prime[49]   = 16'h00E9;
rom_prime[50]   = 16'h00EF;
rom_prime[51]   = 16'h00F1;
rom_prime[52]   = 16'h00FB;
rom_prime[53]   = 16'h0101;
rom_prime[54]   = 16'h0107;
rom_prime[55]   = 16'h010D;
rom_prime[56]   = 16'h010F;
rom_prime[57]   = 16'h0115;
rom_prime[58]   = 16'h0119;
rom_prime[59]   = 16'h011B;
rom_prime[60]   = 16'h0125;
rom_prime[61]   = 16'h0133;
rom_prime[62]   = 16'h0137;
rom_prime[63]   = 16'h0139;
rom_prime[64]   = 16'h013D;
rom_prime[65]   = 16'h014B;
rom_prime[66]   = 16'h0151;
rom_prime[67]   = 16'h015B;
rom_prime[68]   = 16'h015D;
rom_prime[69]   = 16'h0161;
rom_prime[70]   = 16'h0167;
rom_prime[71]   = 16'h016F;
rom_prime[72]   = 16'h0175;
rom_prime[73]   = 16'h017B;
rom_prime[74]   = 16'h017F;
rom_prime[75]   = 16'h0185;
rom_prime[76]   = 16'h018D;
rom_prime[77]   = 16'h0191;
rom_prime[78]   = 16'h0199;
rom_prime[79]   = 16'h01A3;
rom_prime[80]   = 16'h01A5;
rom_prime[81]   = 16'h01AF;
rom_prime[82]   = 16'h01B1;
rom_prime[83]   = 16'h01B7;
rom_prime[84]   = 16'h01BB;
rom_prime[85]   = 16'h01C1;
rom_prime[86]   = 16'h01C9;
rom_prime[87]   = 16'h01CD;
rom_prime[88]   = 16'h01CF;
rom_prime[89]   = 16'h01D3;
rom_prime[90]   = 16'h01DF;
rom_prime[91]   = 16'h01E7;
rom_prime[92]   = 16'h01EB;
rom_prime[93]   = 16'h01F3;
rom_prime[94]   = 16'h01F7;
rom_prime[95]   = 16'h01FD;
rom_prime[96]   = 16'h0209;
rom_prime[97]   = 16'h020B;
rom_prime[98]   = 16'h021D;
rom_prime[99]   = 16'h0223;
rom_prime[100]  = 16'h022D;
rom_prime[101]  = 16'h0233;
rom_prime[102]  = 16'h0239;
rom_prime[103]  = 16'h023B;
rom_prime[104]  = 16'h0241;
rom_prime[105]  = 16'h024B;
rom_prime[106]  = 16'h0251;
rom_prime[107]  = 16'h0257;
rom_prime[108]  = 16'h0259;
rom_prime[109]  = 16'h025F;
rom_prime[110]  = 16'h0265;
rom_prime[111]  = 16'h0269;
rom_prime[112]  = 16'h026B;
rom_prime[113]  = 16'h0277;
rom_prime[114]  = 16'h0281;
rom_prime[115]  = 16'h0283;
rom_prime[116]  = 16'h0287;
rom_prime[117]  = 16'h028D;
rom_prime[118]  = 16'h0293;
rom_prime[119]  = 16'h0295;
rom_prime[120]  = 16'h02A1;
rom_prime[121]  = 16'h02A5;
rom_prime[122]  = 16'h02AB;
rom_prime[123]  = 16'h02B3;
rom_prime[124]  = 16'h02BD;
rom_prime[125]  = 16'h02C5;
rom_prime[126]  = 16'h02CF;
rom_prime[127]  = 16'h02D7;
rom_prime[128]  = 16'h02DD;
rom_prime[129]  = 16'h02E3;
rom_prime[130]  = 16'h02E7;
rom_prime[131]  = 16'h02EF;
rom_prime[132]  = 16'h02F5;
rom_prime[133]  = 16'h02F9;
rom_prime[134]  = 16'h0301;
rom_prime[135]  = 16'h0305;
rom_prime[136]  = 16'h0313;
rom_prime[137]  = 16'h031D;
rom_prime[138]  = 16'h0329;
rom_prime[139]  = 16'h032B;
rom_prime[140]  = 16'h0335;
rom_prime[141]  = 16'h0337;
rom_prime[142]  = 16'h033B;
rom_prime[143]  = 16'h033D;
rom_prime[144]  = 16'h0347;
rom_prime[145]  = 16'h0355;
rom_prime[146]  = 16'h0359;
rom_prime[147]  = 16'h035B;
rom_prime[148]  = 16'h035F;
rom_prime[149]  = 16'h036D;
rom_prime[150]  = 16'h0371;
rom_prime[151]  = 16'h0373;
rom_prime[152]  = 16'h0377;
rom_prime[153]  = 16'h038B;
rom_prime[154]  = 16'h038F;
rom_prime[155]  = 16'h0397;
rom_prime[156]  = 16'h03A1;
rom_prime[157]  = 16'h03A9;
rom_prime[158]  = 16'h03AD;
rom_prime[159]  = 16'h03B3;
rom_prime[160]  = 16'h03B9;
rom_prime[161]  = 16'h03C7;
rom_prime[162]  = 16'h03CB;
rom_prime[163]  = 16'h03D1;
rom_prime[164]  = 16'h03D7;
rom_prime[165]  = 16'h03DF;
rom_prime[166]  = 16'h03E5;
rom_prime[167]  = 16'h03F1;
rom_prime[168]  = 16'h03F5;
rom_prime[169]  = 16'h03FB;
rom_prime[170]  = 16'h03FD;
rom_prime[171]  = 16'h0407;
rom_prime[172]  = 16'h0409;
rom_prime[173]  = 16'h040F;
rom_prime[174]  = 16'h0419;
rom_prime[175]  = 16'h041B;
rom_prime[176]  = 16'h0425;
rom_prime[177]  = 16'h0427;
rom_prime[178]  = 16'h042D;
rom_prime[179]  = 16'h043F;
rom_prime[180]  = 16'h0443;
rom_prime[181]  = 16'h0445;
rom_prime[182]  = 16'h0449;
rom_prime[183]  = 16'h044F;
rom_prime[184]  = 16'h0455;
rom_prime[185]  = 16'h045D;
rom_prime[186]  = 16'h0463;
rom_prime[187]  = 16'h0469;
rom_prime[188]  = 16'h047F;
rom_prime[189]  = 16'h0481;
rom_prime[190]  = 16'h048B;
rom_prime[191]  = 16'h0493;
rom_prime[192]  = 16'h049D;
rom_prime[193]  = 16'h04A3;
rom_prime[194]  = 16'h04A9;
rom_prime[195]  = 16'h04B1;
rom_prime[196]  = 16'h04BD;
rom_prime[197]  = 16'h04C1;
rom_prime[198]  = 16'h04C7;
rom_prime[199]  = 16'h04CD;
rom_prime[200]  = 16'h04CF;
rom_prime[201]  = 16'h04D5;
rom_prime[202]  = 16'h04E1;
rom_prime[203]  = 16'h04EB;
rom_prime[204]  = 16'h04FD;
rom_prime[205]  = 16'h04FF;
rom_prime[206]  = 16'h0503;
rom_prime[207]  = 16'h0509;
rom_prime[208]  = 16'h050B;
rom_prime[209]  = 16'h0511;
rom_prime[210]  = 16'h0515;
rom_prime[211]  = 16'h0517;
rom_prime[212]  = 16'h051B;
rom_prime[213]  = 16'h0527;
rom_prime[214]  = 16'h0529;
rom_prime[215]  = 16'h052F;
rom_prime[216]  = 16'h0551;
rom_prime[217]  = 16'h0557;
rom_prime[218]  = 16'h055D;
rom_prime[219]  = 16'h0565;
rom_prime[220]  = 16'h0577;
rom_prime[221]  = 16'h0581;
rom_prime[222]  = 16'h058F;
rom_prime[223]  = 16'h0593;
rom_prime[224]  = 16'h0595;
rom_prime[225]  = 16'h0599;
rom_prime[226]  = 16'h059F;
rom_prime[227]  = 16'h05A7;
rom_prime[228]  = 16'h05AB;
rom_prime[229]  = 16'h05AD;
rom_prime[230]  = 16'h05B3;
rom_prime[231]  = 16'h05BF;
rom_prime[232]  = 16'h05C9;
rom_prime[233]  = 16'h05CB;
rom_prime[234]  = 16'h05CF;
rom_prime[235]  = 16'h05D1;
rom_prime[236]  = 16'h05D5;
rom_prime[237]  = 16'h05DB;
rom_prime[238]  = 16'h05E7;
rom_prime[239]  = 16'h05F3;
rom_prime[240]  = 16'h05FB;
rom_prime[241]  = 16'h0607;
rom_prime[242]  = 16'h060D;
rom_prime[243]  = 16'h0611;
rom_prime[244]  = 16'h0617;
rom_prime[245]  = 16'h061F;
rom_prime[246]  = 16'h0623;
rom_prime[247]  = 16'h062B;
rom_prime[248]  = 16'h062F;
rom_prime[249]  = 16'h063D;
rom_prime[250]  = 16'h0641;
rom_prime[251]  = 16'h0647;
rom_prime[252]  = 16'h0649;
rom_prime[253]  = 16'h064D;
rom_prime[254]  = 16'h0653;
rom_prime[255]  = 16'h0655;
rom_prime[256]  = 16'h065B;
rom_prime[257]  = 16'h0665;
rom_prime[258]  = 16'h0679;
rom_prime[259]  = 16'h067F;
rom_prime[260]  = 16'h0683;
rom_prime[261]  = 16'h0685;
rom_prime[262]  = 16'h069D;
rom_prime[263]  = 16'h06A1;
rom_prime[264]  = 16'h06A3;
rom_prime[265]  = 16'h06AD;
rom_prime[266]  = 16'h06B9;
rom_prime[267]  = 16'h06BB;
rom_prime[268]  = 16'h06C5;
rom_prime[269]  = 16'h06CD;
rom_prime[270]  = 16'h06D3;
rom_prime[271]  = 16'h06D9;
rom_prime[272]  = 16'h06DF;
rom_prime[273]  = 16'h06F1;
rom_prime[274]  = 16'h06F7;
rom_prime[275]  = 16'h06FB;
rom_prime[276]  = 16'h06FD;
rom_prime[277]  = 16'h0709;
rom_prime[278]  = 16'h0713;
rom_prime[279]  = 16'h071F;
rom_prime[280]  = 16'h0727;
rom_prime[281]  = 16'h0737;
rom_prime[282]  = 16'h0745;
rom_prime[283]  = 16'h074B;
rom_prime[284]  = 16'h074F;
rom_prime[285]  = 16'h0751;
rom_prime[286]  = 16'h0755;
rom_prime[287]  = 16'h0757;
rom_prime[288]  = 16'h0761;
rom_prime[289]  = 16'h076D;
rom_prime[290]  = 16'h0773;
rom_prime[291]  = 16'h0779;
rom_prime[292]  = 16'h078B;
rom_prime[293]  = 16'h078D;
rom_prime[294]  = 16'h079D;
rom_prime[295]  = 16'h079F;
rom_prime[296]  = 16'h07B5;
rom_prime[297]  = 16'h07BB;
rom_prime[298]  = 16'h07C3;
rom_prime[299]  = 16'h07C9;
rom_prime[300]  = 16'h07CD;
rom_prime[301]  = 16'h07CF;
rom_prime[302]  = 16'h07D3;
rom_prime[303]  = 16'h07DB;
rom_prime[304]  = 16'h07E1;
rom_prime[305]  = 16'h07EB;
rom_prime[306]  = 16'h07ED;
rom_prime[307]  = 16'h07F7;
rom_prime[308]  = 16'h0805;
rom_prime[309]  = 16'h080F;
rom_prime[310]  = 16'h0815;
rom_prime[311]  = 16'h0821;
rom_prime[312]  = 16'h0823;
rom_prime[313]  = 16'h0827;
rom_prime[314]  = 16'h0829;
rom_prime[315]  = 16'h0833;
rom_prime[316]  = 16'h083F;
rom_prime[317]  = 16'h0841;
rom_prime[318]  = 16'h0851;
rom_prime[319]  = 16'h0853;
rom_prime[320]  = 16'h0859;
rom_prime[321]  = 16'h085D;
rom_prime[322]  = 16'h085F;
rom_prime[323]  = 16'h0869;
rom_prime[324]  = 16'h0871;
rom_prime[325]  = 16'h0883;
rom_prime[326]  = 16'h089B;
rom_prime[327]  = 16'h089F;
rom_prime[328]  = 16'h08A5;
rom_prime[329]  = 16'h08AD;
rom_prime[330]  = 16'h08BD;
rom_prime[331]  = 16'h08BF;
rom_prime[332]  = 16'h08C3;
rom_prime[333]  = 16'h08CB;
rom_prime[334]  = 16'h08DB;
rom_prime[335]  = 16'h08DD;
rom_prime[336]  = 16'h08E1;
rom_prime[337]  = 16'h08E9;
rom_prime[338]  = 16'h08EF;
rom_prime[339]  = 16'h08F5;
rom_prime[340]  = 16'h08F9;
rom_prime[341]  = 16'h0905;
rom_prime[342]  = 16'h0907;
rom_prime[343]  = 16'h091D;
rom_prime[344]  = 16'h0923;
rom_prime[345]  = 16'h0925;
rom_prime[346]  = 16'h092B;
rom_prime[347]  = 16'h092F;
rom_prime[348]  = 16'h0935;
rom_prime[349]  = 16'h0943;
rom_prime[350]  = 16'h0949;
rom_prime[351]  = 16'h094D;
rom_prime[352]  = 16'h094F;
rom_prime[353]  = 16'h0955;
rom_prime[354]  = 16'h0959;
rom_prime[355]  = 16'h095F;
rom_prime[356]  = 16'h096B;
rom_prime[357]  = 16'h0971;
rom_prime[358]  = 16'h0977;
rom_prime[359]  = 16'h0985;
rom_prime[360]  = 16'h0989;
rom_prime[361]  = 16'h098F;
rom_prime[362]  = 16'h099B;
rom_prime[363]  = 16'h09A3;
rom_prime[364]  = 16'h09A9;
rom_prime[365]  = 16'h09AD;
rom_prime[366]  = 16'h09C7;
rom_prime[367]  = 16'h09D9;
rom_prime[368]  = 16'h09E3;
rom_prime[369]  = 16'h09EB;
rom_prime[370]  = 16'h09EF;
rom_prime[371]  = 16'h09F5;
rom_prime[372]  = 16'h09F7;
rom_prime[373]  = 16'h09FD;
rom_prime[374]  = 16'h0A13;
rom_prime[375]  = 16'h0A1F;
rom_prime[376]  = 16'h0A21;
rom_prime[377]  = 16'h0A31;
rom_prime[378]  = 16'h0A39;
rom_prime[379]  = 16'h0A3D;
rom_prime[380]  = 16'h0A49;
rom_prime[381]  = 16'h0A57;
rom_prime[382]  = 16'h0A61;
rom_prime[383]  = 16'h0A63;
rom_prime[384]  = 16'h0A67;
rom_prime[385]  = 16'h0A6F;
rom_prime[386]  = 16'h0A75;
rom_prime[387]  = 16'h0A7B;
rom_prime[388]  = 16'h0A7F;
rom_prime[389]  = 16'h0A81;
rom_prime[390]  = 16'h0A85;
rom_prime[391]  = 16'h0A8B;
rom_prime[392]  = 16'h0A93;
rom_prime[393]  = 16'h0A97;
rom_prime[394]  = 16'h0A99;
rom_prime[395]  = 16'h0A9F;
rom_prime[396]  = 16'h0AA9;
rom_prime[397]  = 16'h0AAB;
rom_prime[398]  = 16'h0AB5;
rom_prime[399]  = 16'h0ABD;
rom_prime[400]  = 16'h0AC1;
rom_prime[401]  = 16'h0ACF;
rom_prime[402]  = 16'h0AD9;
rom_prime[403]  = 16'h0AE5;
rom_prime[404]  = 16'h0AE7;
rom_prime[405]  = 16'h0AED;
rom_prime[406]  = 16'h0AF1;
rom_prime[407]  = 16'h0AF3;
rom_prime[408]  = 16'h0B03;
rom_prime[409]  = 16'h0B11;
rom_prime[410]  = 16'h0B15;
rom_prime[411]  = 16'h0B1B;
rom_prime[412]  = 16'h0B23;
rom_prime[413]  = 16'h0B29;
rom_prime[414]  = 16'h0B2D;
rom_prime[415]  = 16'h0B3F;
rom_prime[416]  = 16'h0B47;
rom_prime[417]  = 16'h0B51;
rom_prime[418]  = 16'h0B57;
rom_prime[419]  = 16'h0B5D;
rom_prime[420]  = 16'h0B65;
rom_prime[421]  = 16'h0B6F;
rom_prime[422]  = 16'h0B7B;
rom_prime[423]  = 16'h0B89;
rom_prime[424]  = 16'h0B8D;
rom_prime[425]  = 16'h0B93;
rom_prime[426]  = 16'h0B99;
rom_prime[427]  = 16'h0B9B;
rom_prime[428]  = 16'h0BB7;
rom_prime[429]  = 16'h0BB9;
rom_prime[430]  = 16'h0BC3;
rom_prime[431]  = 16'h0BCB;
rom_prime[432]  = 16'h0BCF;
rom_prime[433]  = 16'h0BDD;
rom_prime[434]  = 16'h0BE1;
rom_prime[435]  = 16'h0BE9;
rom_prime[436]  = 16'h0BF5;
rom_prime[437]  = 16'h0BFB;
rom_prime[438]  = 16'h0C07;
rom_prime[439]  = 16'h0C0B;
rom_prime[440]  = 16'h0C11;
rom_prime[441]  = 16'h0C25;
rom_prime[442]  = 16'h0C2F;
rom_prime[443]  = 16'h0C31;
rom_prime[444]  = 16'h0C41;
rom_prime[445]  = 16'h0C5B;
rom_prime[446]  = 16'h0C5F;
rom_prime[447]  = 16'h0C61;
rom_prime[448]  = 16'h0C6D;
rom_prime[449]  = 16'h0C73;
rom_prime[450]  = 16'h0C77;
rom_prime[451]  = 16'h0C83;
rom_prime[452]  = 16'h0C89;
rom_prime[453]  = 16'h0C91;
rom_prime[454]  = 16'h0C95;
rom_prime[455]  = 16'h0C9D;
rom_prime[456]  = 16'h0CB3;
rom_prime[457]  = 16'h0CB5;
rom_prime[458]  = 16'h0CB9;
rom_prime[459]  = 16'h0CBB;
rom_prime[460]  = 16'h0CC7;
rom_prime[461]  = 16'h0CE3;
rom_prime[462]  = 16'h0CE5;
rom_prime[463]  = 16'h0CEB;
rom_prime[464]  = 16'h0CF1;
rom_prime[465]  = 16'h0CF7;
rom_prime[466]  = 16'h0CFB;
rom_prime[467]  = 16'h0D01;
rom_prime[468]  = 16'h0D03;
rom_prime[469]  = 16'h0D0F;
rom_prime[470]  = 16'h0D13;
rom_prime[471]  = 16'h0D1F;
rom_prime[472]  = 16'h0D21;
rom_prime[473]  = 16'h0D2B;
rom_prime[474]  = 16'h0D2D;
rom_prime[475]  = 16'h0D3D;
rom_prime[476]  = 16'h0D3F;
rom_prime[477]  = 16'h0D4F;
rom_prime[478]  = 16'h0D55;
rom_prime[479]  = 16'h0D69;
rom_prime[480]  = 16'h0D79;
rom_prime[481]  = 16'h0D81;
rom_prime[482]  = 16'h0D85;
rom_prime[483]  = 16'h0D87;
rom_prime[484]  = 16'h0D8B;
rom_prime[485]  = 16'h0D8D;
rom_prime[486]  = 16'h0DA3;
rom_prime[487]  = 16'h0DAB;
rom_prime[488]  = 16'h0DB7;
rom_prime[489]  = 16'h0DBD;
rom_prime[490]  = 16'h0DC7;
rom_prime[491]  = 16'h0DC9;
rom_prime[492]  = 16'h0DCD;
rom_prime[493]  = 16'h0DD3;
rom_prime[494]  = 16'h0DD5;
rom_prime[495]  = 16'h0DDB;
rom_prime[496]  = 16'h0DE5;
rom_prime[497]  = 16'h0DE7;
rom_prime[498]  = 16'h0DF3;
rom_prime[499]  = 16'h0DFD;
rom_prime[500]  = 16'h0DFF;
rom_prime[501]  = 16'h0E09;
rom_prime[502]  = 16'h0E17;
rom_prime[503]  = 16'h0E1D;
rom_prime[504]  = 16'h0E21;
rom_prime[505]  = 16'h0E27;
rom_prime[506]  = 16'h0E2F;
rom_prime[507]  = 16'h0E35;
rom_prime[508]  = 16'h0E3B;
rom_prime[509]  = 16'h0E4B;
rom_prime[510]  = 16'h0E57;
rom_prime[511]  = 16'h0E59;
rom_prime[512]  = 16'h0E5D;
rom_prime[513]  = 16'h0E6B;
rom_prime[514]  = 16'h0E71;
rom_prime[515]  = 16'h0E75;
rom_prime[516]  = 16'h0E7D;
rom_prime[517]  = 16'h0E87;
rom_prime[518]  = 16'h0E8F;
rom_prime[519]  = 16'h0E95;
rom_prime[520]  = 16'h0E9B;
rom_prime[521]  = 16'h0EB1;
rom_prime[522]  = 16'h0EB7;
rom_prime[523]  = 16'h0EB9;
rom_prime[524]  = 16'h0EC3;
rom_prime[525]  = 16'h0ED1;
rom_prime[526]  = 16'h0ED5;
rom_prime[527]  = 16'h0EDB;
rom_prime[528]  = 16'h0EED;
rom_prime[529]  = 16'h0EEF;
rom_prime[530]  = 16'h0EF9;
rom_prime[531]  = 16'h0F07;
rom_prime[532]  = 16'h0F0B;
rom_prime[533]  = 16'h0F0D;
rom_prime[534]  = 16'h0F17;
rom_prime[535]  = 16'h0F25;
rom_prime[536]  = 16'h0F29;
rom_prime[537]  = 16'h0F31;
rom_prime[538]  = 16'h0F43;
rom_prime[539]  = 16'h0F47;
rom_prime[540]  = 16'h0F4D;
rom_prime[541]  = 16'h0F4F;
rom_prime[542]  = 16'h0F53;
rom_prime[543]  = 16'h0F59;
rom_prime[544]  = 16'h0F5B;
rom_prime[545]  = 16'h0F67;
rom_prime[546]  = 16'h0F6B;
rom_prime[547]  = 16'h0F7F;
rom_prime[548]  = 16'h0F95;
rom_prime[549]  = 16'h0FA1;
rom_prime[550]  = 16'h0FA3;
rom_prime[551]  = 16'h0FA7;
rom_prime[552]  = 16'h0FAD;
rom_prime[553]  = 16'h0FB3;
rom_prime[554]  = 16'h0FB5;
rom_prime[555]  = 16'h0FBB;
rom_prime[556]  = 16'h0FD1;
rom_prime[557]  = 16'h0FD3;
rom_prime[558]  = 16'h0FD9;
rom_prime[559]  = 16'h0FE9;
rom_prime[560]  = 16'h0FEF;
rom_prime[561]  = 16'h0FFB;
rom_prime[562]  = 16'h0FFD;
rom_prime[563]  = 16'h1003;
rom_prime[564]  = 16'h100F;
rom_prime[565]  = 16'h101F;
rom_prime[566]  = 16'h1021;
rom_prime[567]  = 16'h1025;
rom_prime[568]  = 16'h102B;
rom_prime[569]  = 16'h1039;
rom_prime[570]  = 16'h103D;
rom_prime[571]  = 16'h103F;
rom_prime[572]  = 16'h1051;
rom_prime[573]  = 16'h1069;
rom_prime[574]  = 16'h1073;
rom_prime[575]  = 16'h1079;
rom_prime[576]  = 16'h107B;
rom_prime[577]  = 16'h1085;
rom_prime[578]  = 16'h1087;
rom_prime[579]  = 16'h1091;
rom_prime[580]  = 16'h1093;
rom_prime[581]  = 16'h109D;
rom_prime[582]  = 16'h10A3;
rom_prime[583]  = 16'h10A5;
rom_prime[584]  = 16'h10AF;
rom_prime[585]  = 16'h10B1;
rom_prime[586]  = 16'h10BB;
rom_prime[587]  = 16'h10C1;
rom_prime[588]  = 16'h10C9;
rom_prime[589]  = 16'h10E7;
rom_prime[590]  = 16'h10F1;
rom_prime[591]  = 16'h10F3;
rom_prime[592]  = 16'h10FD;
rom_prime[593]  = 16'h1105;
rom_prime[594]  = 16'h110B;
rom_prime[595]  = 16'h1115;
rom_prime[596]  = 16'h1127;
rom_prime[597]  = 16'h112D;
rom_prime[598]  = 16'h1139;
rom_prime[599]  = 16'h1145;
rom_prime[600]  = 16'h1147;
rom_prime[601]  = 16'h1159;
rom_prime[602]  = 16'h115F;
rom_prime[603]  = 16'h1163;
rom_prime[604]  = 16'h1169;
rom_prime[605]  = 16'h116F;
rom_prime[606]  = 16'h1181;
rom_prime[607]  = 16'h1183;
rom_prime[608]  = 16'h118D;
rom_prime[609]  = 16'h119B;
rom_prime[610]  = 16'h11A1;
rom_prime[611]  = 16'h11A5;
rom_prime[612]  = 16'h11A7;
rom_prime[613]  = 16'h11AB;
rom_prime[614]  = 16'h11C3;
rom_prime[615]  = 16'h11C5;
rom_prime[616]  = 16'h11D1;
rom_prime[617]  = 16'h11D7;
rom_prime[618]  = 16'h11E7;
rom_prime[619]  = 16'h11EF;
rom_prime[620]  = 16'h11F5;
rom_prime[621]  = 16'h11FB;
rom_prime[622]  = 16'h120D;
rom_prime[623]  = 16'h121D;
rom_prime[624]  = 16'h121F;
rom_prime[625]  = 16'h1223;
rom_prime[626]  = 16'h1229;
rom_prime[627]  = 16'h122B;
rom_prime[628]  = 16'h1231;
rom_prime[629]  = 16'h1237;
rom_prime[630]  = 16'h1241;
rom_prime[631]  = 16'h1247;
rom_prime[632]  = 16'h1253;
rom_prime[633]  = 16'h125F;
rom_prime[634]  = 16'h1271;
rom_prime[635]  = 16'h1273;
rom_prime[636]  = 16'h1279;
rom_prime[637]  = 16'h127D;
rom_prime[638]  = 16'h128F;
rom_prime[639]  = 16'h1297;
rom_prime[640]  = 16'h12AF;
rom_prime[641]  = 16'h12B3;
rom_prime[642]  = 16'h12B5;
rom_prime[643]  = 16'h12B9;
rom_prime[644]  = 16'h12BF;
rom_prime[645]  = 16'h12C1;
rom_prime[646]  = 16'h12CD;
rom_prime[647]  = 16'h12D1;
rom_prime[648]  = 16'h12DF;
rom_prime[649]  = 16'h12FD;
rom_prime[650]  = 16'h1307;
rom_prime[651]  = 16'h130D;
rom_prime[652]  = 16'h1319;
rom_prime[653]  = 16'h1327;
rom_prime[654]  = 16'h132D;
rom_prime[655]  = 16'h1337;
rom_prime[656]  = 16'h1343;
rom_prime[657]  = 16'h1345;
rom_prime[658]  = 16'h1349;
rom_prime[659]  = 16'h134F;
rom_prime[660]  = 16'h1357;
rom_prime[661]  = 16'h135D;
rom_prime[662]  = 16'h1367;
rom_prime[663]  = 16'h1369;
rom_prime[664]  = 16'h136D;
rom_prime[665]  = 16'h137B;
rom_prime[666]  = 16'h1381;
rom_prime[667]  = 16'h1387;
rom_prime[668]  = 16'h138B;
rom_prime[669]  = 16'h1391;
rom_prime[670]  = 16'h1393;
rom_prime[671]  = 16'h139D;
rom_prime[672]  = 16'h139F;
rom_prime[673]  = 16'h13AF;
rom_prime[674]  = 16'h13BB;
rom_prime[675]  = 16'h13C3;
rom_prime[676]  = 16'h13D5;
rom_prime[677]  = 16'h13D9;
rom_prime[678]  = 16'h13DF;
rom_prime[679]  = 16'h13EB;
rom_prime[680]  = 16'h13ED;
rom_prime[681]  = 16'h13F3;
rom_prime[682]  = 16'h13F9;
rom_prime[683]  = 16'h13FF;
rom_prime[684]  = 16'h141B;
rom_prime[685]  = 16'h1421;
rom_prime[686]  = 16'h142F;
rom_prime[687]  = 16'h1433;
rom_prime[688]  = 16'h143B;
rom_prime[689]  = 16'h1445;
rom_prime[690]  = 16'h144D;
rom_prime[691]  = 16'h1459;
rom_prime[692]  = 16'h146B;
rom_prime[693]  = 16'h146F;
rom_prime[694]  = 16'h1471;
rom_prime[695]  = 16'h1475;
rom_prime[696]  = 16'h148D;
rom_prime[697]  = 16'h1499;
rom_prime[698]  = 16'h149F;
rom_prime[699]  = 16'h14A1;
rom_prime[700]  = 16'h14B1;
rom_prime[701]  = 16'h14B7;
rom_prime[702]  = 16'h14BD;
rom_prime[703]  = 16'h14CB;
rom_prime[704]  = 16'h14D5;
rom_prime[705]  = 16'h14E3;
rom_prime[706]  = 16'h14E7;
rom_prime[707]  = 16'h1505;
rom_prime[708]  = 16'h150B;
rom_prime[709]  = 16'h1511;
rom_prime[710]  = 16'h1517;
rom_prime[711]  = 16'h151F;
rom_prime[712]  = 16'h1525;
rom_prime[713]  = 16'h1529;
rom_prime[714]  = 16'h152B;
rom_prime[715]  = 16'h1537;
rom_prime[716]  = 16'h153D;
rom_prime[717]  = 16'h1541;
rom_prime[718]  = 16'h1543;
rom_prime[719]  = 16'h1549;
rom_prime[720]  = 16'h155F;
rom_prime[721]  = 16'h1565;
rom_prime[722]  = 16'h1567;
rom_prime[723]  = 16'h156B;
rom_prime[724]  = 16'h157D;
rom_prime[725]  = 16'h157F;
rom_prime[726]  = 16'h1583;
rom_prime[727]  = 16'h158F;
rom_prime[728]  = 16'h1591;
rom_prime[729]  = 16'h1597;
rom_prime[730]  = 16'h159B;
rom_prime[731]  = 16'h15B5;
rom_prime[732]  = 16'h15BB;
rom_prime[733]  = 16'h15C1;
rom_prime[734]  = 16'h15C5;
rom_prime[735]  = 16'h15CD;
rom_prime[736]  = 16'h15D7;
rom_prime[737]  = 16'h15F7;
rom_prime[738]  = 16'h1607;
rom_prime[739]  = 16'h1609;
rom_prime[740]  = 16'h160F;
rom_prime[741]  = 16'h1613;
rom_prime[742]  = 16'h1615;
rom_prime[743]  = 16'h1619;
rom_prime[744]  = 16'h161B;
rom_prime[745]  = 16'h1625;
rom_prime[746]  = 16'h1633;
rom_prime[747]  = 16'h1639;
rom_prime[748]  = 16'h163D;
rom_prime[749]  = 16'h1645;
rom_prime[750]  = 16'h164F;
rom_prime[751]  = 16'h1655;
rom_prime[752]  = 16'h1669;
rom_prime[753]  = 16'h166D;
rom_prime[754]  = 16'h166F;
rom_prime[755]  = 16'h1675;
rom_prime[756]  = 16'h1693;
rom_prime[757]  = 16'h1697;
rom_prime[758]  = 16'h169F;
rom_prime[759]  = 16'h16A9;
rom_prime[760]  = 16'h16AF;
rom_prime[761]  = 16'h16B5;
rom_prime[762]  = 16'h16BD;
rom_prime[763]  = 16'h16C3;
rom_prime[764]  = 16'h16CF;
rom_prime[765]  = 16'h16D3;
rom_prime[766]  = 16'h16D9;
rom_prime[767]  = 16'h16DB;
rom_prime[768]  = 16'h16E1;
rom_prime[769]  = 16'h16E5;
rom_prime[770]  = 16'h16EB;
rom_prime[771]  = 16'h16ED;
rom_prime[772]  = 16'h16F7;
rom_prime[773]  = 16'h16F9;
rom_prime[774]  = 16'h1709;
rom_prime[775]  = 16'h170F;
rom_prime[776]  = 16'h1723;
rom_prime[777]  = 16'h1727;
rom_prime[778]  = 16'h1733;
rom_prime[779]  = 16'h1741;
rom_prime[780]  = 16'h175D;
rom_prime[781]  = 16'h1763;
rom_prime[782]  = 16'h1777;
rom_prime[783]  = 16'h177B;
rom_prime[784]  = 16'h178D;
rom_prime[785]  = 16'h1795;
rom_prime[786]  = 16'h179B;
rom_prime[787]  = 16'h179F;
rom_prime[788]  = 16'h17A5;
rom_prime[789]  = 16'h17B3;
rom_prime[790]  = 16'h17B9;
rom_prime[791]  = 16'h17BF;
rom_prime[792]  = 16'h17C9;
rom_prime[793]  = 16'h17CB;
rom_prime[794]  = 16'h17D5;
rom_prime[795]  = 16'h17E1;
rom_prime[796]  = 16'h17E9;
rom_prime[797]  = 16'h17F3;
rom_prime[798]  = 16'h17F5;
rom_prime[799]  = 16'h17FF;
rom_prime[800]  = 16'h1807;
rom_prime[801]  = 16'h1813;
rom_prime[802]  = 16'h181D;
rom_prime[803]  = 16'h1835;
rom_prime[804]  = 16'h1837;
rom_prime[805]  = 16'h183B;
rom_prime[806]  = 16'h1843;
rom_prime[807]  = 16'h1849;
rom_prime[808]  = 16'h184D;
rom_prime[809]  = 16'h1855;
rom_prime[810]  = 16'h1867;
rom_prime[811]  = 16'h1871;
rom_prime[812]  = 16'h1877;
rom_prime[813]  = 16'h187D;
rom_prime[814]  = 16'h187F;
rom_prime[815]  = 16'h1885;
rom_prime[816]  = 16'h188F;
rom_prime[817]  = 16'h189B;
rom_prime[818]  = 16'h189D;
rom_prime[819]  = 16'h18A7;
rom_prime[820]  = 16'h18AD;
rom_prime[821]  = 16'h18B3;
rom_prime[822]  = 16'h18B9;
rom_prime[823]  = 16'h18C1;
rom_prime[824]  = 16'h18C7;
rom_prime[825]  = 16'h18D1;
rom_prime[826]  = 16'h18D7;
rom_prime[827]  = 16'h18D9;
rom_prime[828]  = 16'h18DF;
rom_prime[829]  = 16'h18E5;
rom_prime[830]  = 16'h18EB;
rom_prime[831]  = 16'h18F5;
rom_prime[832]  = 16'h18FD;
rom_prime[833]  = 16'h1915;
rom_prime[834]  = 16'h191B;
rom_prime[835]  = 16'h1931;
rom_prime[836]  = 16'h1933;
rom_prime[837]  = 16'h1945;
rom_prime[838]  = 16'h1949;
rom_prime[839]  = 16'h1951;
rom_prime[840]  = 16'h195B;
rom_prime[841]  = 16'h1979;
rom_prime[842]  = 16'h1981;
rom_prime[843]  = 16'h1993;
rom_prime[844]  = 16'h1997;
rom_prime[845]  = 16'h1999;
rom_prime[846]  = 16'h19A3;
rom_prime[847]  = 16'h19A9;
rom_prime[848]  = 16'h19AB;
rom_prime[849]  = 16'h19B1;
rom_prime[850]  = 16'h19B5;
rom_prime[851]  = 16'h19C7;
rom_prime[852]  = 16'h19CF;
rom_prime[853]  = 16'h19DB;
rom_prime[854]  = 16'h19ED;
rom_prime[855]  = 16'h19FD;
rom_prime[856]  = 16'h1A03;
rom_prime[857]  = 16'h1A05;
rom_prime[858]  = 16'h1A11;
rom_prime[859]  = 16'h1A17;
rom_prime[860]  = 16'h1A21;
rom_prime[861]  = 16'h1A23;
rom_prime[862]  = 16'h1A2D;
rom_prime[863]  = 16'h1A2F;
rom_prime[864]  = 16'h1A35;
rom_prime[865]  = 16'h1A3F;
rom_prime[866]  = 16'h1A4D;
rom_prime[867]  = 16'h1A51;
rom_prime[868]  = 16'h1A69;
rom_prime[869]  = 16'h1A6B;
rom_prime[870]  = 16'h1A7B;
rom_prime[871]  = 16'h1A7D;
rom_prime[872]  = 16'h1A87;
rom_prime[873]  = 16'h1A89;
rom_prime[874]  = 16'h1A93;
rom_prime[875]  = 16'h1AA7;
rom_prime[876]  = 16'h1AAB;
rom_prime[877]  = 16'h1AAD;
rom_prime[878]  = 16'h1AB1;
rom_prime[879]  = 16'h1AB9;
rom_prime[880]  = 16'h1AC9;
rom_prime[881]  = 16'h1ACF;
rom_prime[882]  = 16'h1AD5;
rom_prime[883]  = 16'h1AD7;
rom_prime[884]  = 16'h1AE3;
rom_prime[885]  = 16'h1AF3;
rom_prime[886]  = 16'h1AFB;
rom_prime[887]  = 16'h1AFF;
rom_prime[888]  = 16'h1B05;
rom_prime[889]  = 16'h1B23;
rom_prime[890]  = 16'h1B25;
rom_prime[891]  = 16'h1B2F;
rom_prime[892]  = 16'h1B31;
rom_prime[893]  = 16'h1B37;
rom_prime[894]  = 16'h1B3B;
rom_prime[895]  = 16'h1B41;
rom_prime[896]  = 16'h1B47;
rom_prime[897]  = 16'h1B4F;
rom_prime[898]  = 16'h1B55;
rom_prime[899]  = 16'h1B59;
rom_prime[900]  = 16'h1B65;
rom_prime[901]  = 16'h1B6B;
rom_prime[902]  = 16'h1B73;
rom_prime[903]  = 16'h1B7F;
rom_prime[904]  = 16'h1B83;
rom_prime[905]  = 16'h1B91;
rom_prime[906]  = 16'h1B9D;
rom_prime[907]  = 16'h1BA7;
rom_prime[908]  = 16'h1BBF;
rom_prime[909]  = 16'h1BC5;
rom_prime[910]  = 16'h1BD1;
rom_prime[911]  = 16'h1BD7;
rom_prime[912]  = 16'h1BD9;
rom_prime[913]  = 16'h1BEF;
rom_prime[914]  = 16'h1BF7;
rom_prime[915]  = 16'h1C09;
rom_prime[916]  = 16'h1C13;
rom_prime[917]  = 16'h1C19;
rom_prime[918]  = 16'h1C27;
rom_prime[919]  = 16'h1C2B;
rom_prime[920]  = 16'h1C2D;
rom_prime[921]  = 16'h1C33;
rom_prime[922]  = 16'h1C3D;
rom_prime[923]  = 16'h1C45;
rom_prime[924]  = 16'h1C4B;
rom_prime[925]  = 16'h1C4F;
rom_prime[926]  = 16'h1C55;
rom_prime[927]  = 16'h1C73;
rom_prime[928]  = 16'h1C81;
rom_prime[929]  = 16'h1C8B;
rom_prime[930]  = 16'h1C8D;
rom_prime[931]  = 16'h1C99;
rom_prime[932]  = 16'h1CA3;
rom_prime[933]  = 16'h1CA5;
rom_prime[934]  = 16'h1CB5;
rom_prime[935]  = 16'h1CB7;
rom_prime[936]  = 16'h1CC9;
rom_prime[937]  = 16'h1CE1;
rom_prime[938]  = 16'h1CF3;
rom_prime[939]  = 16'h1CF9;
rom_prime[940]  = 16'h1D09;
rom_prime[941]  = 16'h1D1B;
rom_prime[942]  = 16'h1D21;
rom_prime[943]  = 16'h1D23;
rom_prime[944]  = 16'h1D35;
rom_prime[945]  = 16'h1D39;
rom_prime[946]  = 16'h1D3F;
rom_prime[947]  = 16'h1D41;
rom_prime[948]  = 16'h1D4B;
rom_prime[949]  = 16'h1D53;
rom_prime[950]  = 16'h1D5D;
rom_prime[951]  = 16'h1D63;
rom_prime[952]  = 16'h1D69;
rom_prime[953]  = 16'h1D71;
rom_prime[954]  = 16'h1D75;
rom_prime[955]  = 16'h1D7B;
rom_prime[956]  = 16'h1D7D;
rom_prime[957]  = 16'h1D87;
rom_prime[958]  = 16'h1D89;
rom_prime[959]  = 16'h1D95;
rom_prime[960]  = 16'h1D99;
rom_prime[961]  = 16'h1D9F;
rom_prime[962]  = 16'h1DA5;
rom_prime[963]  = 16'h1DA7;
rom_prime[964]  = 16'h1DB3;
rom_prime[965]  = 16'h1DB7;
rom_prime[966]  = 16'h1DC5;
rom_prime[967]  = 16'h1DD7;
rom_prime[968]  = 16'h1DDB;
rom_prime[969]  = 16'h1DE1;
rom_prime[970]  = 16'h1DF5;
rom_prime[971]  = 16'h1DF9;
rom_prime[972]  = 16'h1E01;
rom_prime[973]  = 16'h1E07;
rom_prime[974]  = 16'h1E0B;
rom_prime[975]  = 16'h1E13;
rom_prime[976]  = 16'h1E17;
rom_prime[977]  = 16'h1E25;
rom_prime[978]  = 16'h1E2B;
rom_prime[979]  = 16'h1E2F;
rom_prime[980]  = 16'h1E3D;
rom_prime[981]  = 16'h1E49;
rom_prime[982]  = 16'h1E4D;
rom_prime[983]  = 16'h1E4F;
rom_prime[984]  = 16'h1E6D;
rom_prime[985]  = 16'h1E71;
rom_prime[986]  = 16'h1E89;
rom_prime[987]  = 16'h1E8F;
rom_prime[988]  = 16'h1E95;
rom_prime[989]  = 16'h1EA1;
rom_prime[990]  = 16'h1EAD;
rom_prime[991]  = 16'h1EBB;
rom_prime[992]  = 16'h1EC1;
rom_prime[993]  = 16'h1EC5;
rom_prime[994]  = 16'h1EC7;
rom_prime[995]  = 16'h1ECB;
rom_prime[996]  = 16'h1EDD;
rom_prime[997]  = 16'h1EE3;
rom_prime[998]  = 16'h1EEF;
rom_prime[999]  = 16'h1EF7;
rom_prime[1000] = 16'h1EFD;
rom_prime[1001] = 16'h1F01;
rom_prime[1002] = 16'h1F0D;
rom_prime[1003] = 16'h1F0F;
rom_prime[1004] = 16'h1F1B;
rom_prime[1005] = 16'h1F39;
rom_prime[1006] = 16'h1F49;
rom_prime[1007] = 16'h1F4B;
rom_prime[1008] = 16'h1F51;
rom_prime[1009] = 16'h1F67;
rom_prime[1010] = 16'h1F75;
rom_prime[1011] = 16'h1F7B;
rom_prime[1012] = 16'h1F85;
rom_prime[1013] = 16'h1F91;
rom_prime[1014] = 16'h1F97;
rom_prime[1015] = 16'h1F99;
rom_prime[1016] = 16'h1F9D;
rom_prime[1017] = 16'h1FA5;
rom_prime[1018] = 16'h1FAF;
rom_prime[1019] = 16'h1FB5;
rom_prime[1020] = 16'h1FBB;
rom_prime[1021] = 16'h1FD3;
rom_prime[1022] = 16'h1FE1;
rom_prime[1023] = 16'h1FE7;
rom_prime[1024] = 16'h1FEB;
rom_prime[1025] = 16'h1FF3;
rom_prime[1026] = 16'h1FFF;
rom_prime[1027] = 16'h2011;
rom_prime[1028] = 16'h201B;
rom_prime[1029] = 16'h201D;
rom_prime[1030] = 16'h2027;
rom_prime[1031] = 16'h2029;
rom_prime[1032] = 16'h202D;
rom_prime[1033] = 16'h2033;
rom_prime[1034] = 16'h2047;
rom_prime[1035] = 16'h204D;
rom_prime[1036] = 16'h2051;
rom_prime[1037] = 16'h205F;
rom_prime[1038] = 16'h2063;
rom_prime[1039] = 16'h2065;
rom_prime[1040] = 16'h2069;
rom_prime[1041] = 16'h2077;
rom_prime[1042] = 16'h207D;
rom_prime[1043] = 16'h2089;
rom_prime[1044] = 16'h20A1;
rom_prime[1045] = 16'h20AB;
rom_prime[1046] = 16'h20B1;
rom_prime[1047] = 16'h20B9;
rom_prime[1048] = 16'h20C3;
rom_prime[1049] = 16'h20C5;
rom_prime[1050] = 16'h20E3;
rom_prime[1051] = 16'h20E7;
rom_prime[1052] = 16'h20ED;
rom_prime[1053] = 16'h20EF;
rom_prime[1054] = 16'h20FB;
rom_prime[1055] = 16'h20FF;
rom_prime[1056] = 16'h210D;
rom_prime[1057] = 16'h2113;
rom_prime[1058] = 16'h2135;
rom_prime[1059] = 16'h2141;
rom_prime[1060] = 16'h2149;
rom_prime[1061] = 16'h214F;
rom_prime[1062] = 16'h2159;
rom_prime[1063] = 16'h215B;
rom_prime[1064] = 16'h215F;
rom_prime[1065] = 16'h2173;
rom_prime[1066] = 16'h217D;
rom_prime[1067] = 16'h2185;
rom_prime[1068] = 16'h2195;
rom_prime[1069] = 16'h2197;
rom_prime[1070] = 16'h21A1;
rom_prime[1071] = 16'h21AF;
rom_prime[1072] = 16'h21B3;
rom_prime[1073] = 16'h21B5;
rom_prime[1074] = 16'h21C1;
rom_prime[1075] = 16'h21C7;
rom_prime[1076] = 16'h21D7;
rom_prime[1077] = 16'h21DD;
rom_prime[1078] = 16'h21E5;
rom_prime[1079] = 16'h21E9;
rom_prime[1080] = 16'h21F1;
rom_prime[1081] = 16'h21F5;
rom_prime[1082] = 16'h21FB;
rom_prime[1083] = 16'h2203;
rom_prime[1084] = 16'h2209;
rom_prime[1085] = 16'h220F;
rom_prime[1086] = 16'h221B;
rom_prime[1087] = 16'h2221;
rom_prime[1088] = 16'h2225;
rom_prime[1089] = 16'h222B;
rom_prime[1090] = 16'h2231;
rom_prime[1091] = 16'h2239;
rom_prime[1092] = 16'h224B;
rom_prime[1093] = 16'h224F;
rom_prime[1094] = 16'h2263;
rom_prime[1095] = 16'h2267;
rom_prime[1096] = 16'h2273;
rom_prime[1097] = 16'h2275;
rom_prime[1098] = 16'h227F;
rom_prime[1099] = 16'h2285;
rom_prime[1100] = 16'h2287;
rom_prime[1101] = 16'h2291;
rom_prime[1102] = 16'h229D;
rom_prime[1103] = 16'h229F;
rom_prime[1104] = 16'h22A3;
rom_prime[1105] = 16'h22B7;
rom_prime[1106] = 16'h22BD;
rom_prime[1107] = 16'h22DB;
rom_prime[1108] = 16'h22E1;
rom_prime[1109] = 16'h22E5;
rom_prime[1110] = 16'h22ED;
rom_prime[1111] = 16'h22F7;
rom_prime[1112] = 16'h2303;
rom_prime[1113] = 16'h2309;
rom_prime[1114] = 16'h230B;
rom_prime[1115] = 16'h2327;
rom_prime[1116] = 16'h2329;
rom_prime[1117] = 16'h232F;
rom_prime[1118] = 16'h2333;
rom_prime[1119] = 16'h2335;
rom_prime[1120] = 16'h2345;
rom_prime[1121] = 16'h2351;
rom_prime[1122] = 16'h2353;
rom_prime[1123] = 16'h2359;
rom_prime[1124] = 16'h2363;
rom_prime[1125] = 16'h236B;
rom_prime[1126] = 16'h2383;
rom_prime[1127] = 16'h238F;
rom_prime[1128] = 16'h2395;
rom_prime[1129] = 16'h23A7;
rom_prime[1130] = 16'h23AD;
rom_prime[1131] = 16'h23B1;
rom_prime[1132] = 16'h23BF;
rom_prime[1133] = 16'h23C5;
rom_prime[1134] = 16'h23C9;
rom_prime[1135] = 16'h23D5;
rom_prime[1136] = 16'h23DD;
rom_prime[1137] = 16'h23E3;
rom_prime[1138] = 16'h23EF;
rom_prime[1139] = 16'h23F3;
rom_prime[1140] = 16'h23F9;
rom_prime[1141] = 16'h2405;
rom_prime[1142] = 16'h240B;
rom_prime[1143] = 16'h2417;
rom_prime[1144] = 16'h2419;
rom_prime[1145] = 16'h2429;
rom_prime[1146] = 16'h243D;
rom_prime[1147] = 16'h2441;
rom_prime[1148] = 16'h2443;
rom_prime[1149] = 16'h244D;
rom_prime[1150] = 16'h245F;
rom_prime[1151] = 16'h2467;
rom_prime[1152] = 16'h246B;
rom_prime[1153] = 16'h2479;
rom_prime[1154] = 16'h247D;
rom_prime[1155] = 16'h247F;
rom_prime[1156] = 16'h2485;
rom_prime[1157] = 16'h249B;
rom_prime[1158] = 16'h24A1;
rom_prime[1159] = 16'h24AF;
rom_prime[1160] = 16'h24B5;
rom_prime[1161] = 16'h24BB;
rom_prime[1162] = 16'h24C5;
rom_prime[1163] = 16'h24CB;
rom_prime[1164] = 16'h24CD;
rom_prime[1165] = 16'h24D7;
rom_prime[1166] = 16'h24D9;
rom_prime[1167] = 16'h24DD;
rom_prime[1168] = 16'h24DF;
rom_prime[1169] = 16'h24F5;
rom_prime[1170] = 16'h24F7;
rom_prime[1171] = 16'h24FB;
rom_prime[1172] = 16'h2501;
rom_prime[1173] = 16'h2507;
rom_prime[1174] = 16'h2513;
rom_prime[1175] = 16'h2519;
rom_prime[1176] = 16'h2527;
rom_prime[1177] = 16'h2531;
rom_prime[1178] = 16'h253D;
rom_prime[1179] = 16'h2543;
rom_prime[1180] = 16'h254B;
rom_prime[1181] = 16'h254F;
rom_prime[1182] = 16'h2573;
rom_prime[1183] = 16'h2581;
rom_prime[1184] = 16'h258D;
rom_prime[1185] = 16'h2593;
rom_prime[1186] = 16'h2597;
rom_prime[1187] = 16'h259D;
rom_prime[1188] = 16'h259F;
rom_prime[1189] = 16'h25AB;
rom_prime[1190] = 16'h25B1;
rom_prime[1191] = 16'h25BD;
rom_prime[1192] = 16'h25CD;
rom_prime[1193] = 16'h25CF;
rom_prime[1194] = 16'h25D9;
rom_prime[1195] = 16'h25E1;
rom_prime[1196] = 16'h25F7;
rom_prime[1197] = 16'h25F9;
rom_prime[1198] = 16'h2605;
rom_prime[1199] = 16'h260B;
rom_prime[1200] = 16'h260F;
rom_prime[1201] = 16'h2615;
rom_prime[1202] = 16'h2627;
rom_prime[1203] = 16'h2629;
rom_prime[1204] = 16'h2635;
rom_prime[1205] = 16'h263B;
rom_prime[1206] = 16'h263F;
rom_prime[1207] = 16'h264B;
rom_prime[1208] = 16'h2653;
rom_prime[1209] = 16'h2659;
rom_prime[1210] = 16'h2665;
rom_prime[1211] = 16'h2669;
rom_prime[1212] = 16'h266F;
rom_prime[1213] = 16'h267B;
rom_prime[1214] = 16'h2681;
rom_prime[1215] = 16'h2683;
rom_prime[1216] = 16'h268F;
rom_prime[1217] = 16'h269B;
rom_prime[1218] = 16'h269F;
rom_prime[1219] = 16'h26AD;
rom_prime[1220] = 16'h26B3;
rom_prime[1221] = 16'h26C3;
rom_prime[1222] = 16'h26C9;
rom_prime[1223] = 16'h26CB;
rom_prime[1224] = 16'h26D5;
rom_prime[1225] = 16'h26DD;
rom_prime[1226] = 16'h26EF;
rom_prime[1227] = 16'h26F5;
end

/* ============================================================================
 * ROM output
 * ============================================================================*/
always @(posedge CLK) begin
    data_i <= rom_prime[ADDRESS];
end

assign DATA = data_i;

endmodule    //PRIME_ROM